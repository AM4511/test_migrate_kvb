��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*�/ ��Y֫P�.	A��M�bC8�B_)�
�6�+�����l�D$0)σC7W�7�_-��Y`�o�%�B�D�aD����1����b}�"'���,�}G� �:�xt �m%%?/ ������y�����8{7��Ų�2]�O��R�y׻��Rd���r�8���6�0q"����t[�{���W�a��g�^��dk��� �W�j�_R�i�l>gp��UG�Bg�Mk�{!����+�z��0Ҩ�^-oka%�bOH�ObP�����0��Q�@�����[R��;�������3��[�$N�c��r7�M�>pP��I��@hV����
h�8��l�]B��X>Y�C��LcΌ����""f74�R����t�<[]ܵ[ջ`���h��nO$��Co����Gm�N�!��/.�g�"���]g�|Qg+繭~�#��G<F�%/,<4��T���[�\�1%���S�4��X�r�/2�]7��'���D�YN��&��<KW�q�.�c^�I����2�l���(};����#���y�P�b�g��Bz�*,�L�0�P��@ $�]!�� /���c�d��/9�P�����K�Q�?�O'j�v�; �&I�n�p�+��6�����L�ʄiQ�rm��pY�ss<һ�a�%�4<�4��o�u�M��;^��gęT���cfD��!���V�;2�$���rc����B�v~�C����T�����Q?c��kjI�	��c�x8��:�{0�&S��x�tm�0 �t���?���%��k��[�Bt����܆��x�SN�������^.vC�IEmZ���k��D�����-�@:���
���:��<k4���� ����mW�Ωa��/�R? hQl'�?�u:p�30�'�'"�F�?�	�F o��i���K�n��r�S�c?;�M(t�b�܁�����f��}���<�����3�$Hq�&���D��0�Tkc�I�Z�Ĝn�ݯX]J��	l_������=�<�V�_���I�y>	�;l�"Qa��~^��N��e����顉��|�1��`�~p�u8��$�pg5YEcy�������LH�t�,q>�9��ޜ
�������Es���b���(p
g�uYW�\�h���b]�:���Y�p	m��5�����85C?��~�2���A��4H����S6*mGӫ�F���h�(\��� ̛q[�{��/�.WU�H���σ�5܇��x�,i�x���p�ڊ�bLK�C��de�M>B��KN�M��`��++D�<�p#:��n�RW�g�Wh��vI|q������8�Ǉ�bY����~�7�(���euk���D�B_pu�|�$!x�t��6��r�x�vxU>J���ǚ�*���:�b�A�1�B���Il�.%vm[B>xU=
{EH_����h��>�eqC2��Rn�7��7,�b�1�4��qs���g��fSbl��[>g�v6�`<kH�K�a[�)��!��}������/-�D,�a؏�b~� ���:�x~�����ނD� �g�����ʑ��-p5���C%T���&8�=���uV��gHu�W[�C,P��b�N�*k �}[�ڦ��A���o�����+�%;�_�;��<%��x����-H`�8|�`l��¢��d�v!ݥ��	�-�R�Т/�[�^I�G�u	"0̟!�9���f:�G�ڸ8�eЕ��ߐJ�ݓ��shb�8��"�mJc�)�U?��rT�_��=���<ٷ�WDE�Ȳ��2��;j�S�?D@ƚ�eǶv�+*�k2{�����G[Â�^3��]h*��S~0|�D��w��U�,����`q����e����%�s�����X�s��h�ܣ�bLCQ���*����
EJL����h]�6 0��e~H*[�Z��P��f���Н��N0�j��P""��n�7��ۨk�=y���%\�v��d�-$�{���ӯ��u܄H�/=�w��z��4^0�)��/;G	��vٙGD�0%
)fP �����Ȧ�S��/o �:L�)cq�p��V��J��a�"����,eZ���'E@���1�K�u���:�^�ձ���NDv4����MH6J�ex#�-ɷ����1��n*7g�L4�y?�Hj�b!���2��ոd�9e�j|{���ؙ��1{�yv;��n����r�UA�$\!c;}`#��gfo>�5�/�g�X������;1��#���k�Gw��%��U�WV�-stL�P�@���C��'3���c���L�	����z�I��N����*�#>�MY/��Η�4��_&K8�b��>"�6�I��\���0BU��;%�r�:�C��0�޽pF{e�?5�*�?�y]VE�����Th�A�P�������n^x ���^x����h]��4�Z������F^�K�ZK�]�Y^�#*δ[Ef�W�,N�pfݘ�7�
�I�*?��X첃�e��nI��{�c����������/W_:c-�`��WBP�5������-+!��VJ�?�5�t�y(ᄪX5,AC�����&�Lasf����<�s��<��	N�JY�\w�	QǗ
�6Q���ښ��q�4��*�b�b�g�J����x���S/W詳�M��](x����b	$3&��S	�x<]�n�д3Юpl�-�؂a���j�pgO�`Ȗ)1���!�L�䖡�E��s.��y�������;3\���,���_<<Ά�@IF�b|jR�N~��9#�B�CR������9�S5_�=�hJ+��y�N�M!&zX|�{�|VD�ck�O�	��������;-1���gb^U>9'��Eh�'b��������p��x�6�r�2@�ڥ/��\��;K�i�E����d�:��f\�[H��U׹k� �HvޯLr6uZ$o��Cؼ��ۦTd[�<A�<G�Y�BGBR�������c����|	g����N"NH�:[0s�۠8��Ֆ��y��7����z��D��X��ǯ�]�	���&�%8�?�Կvj� ���+Ϯ�pY�=�f'2����@-�i�{8��SW�]�V�J��<D���W��j��؇M�H%����_5c��|�B,��[M���>��%$L���*NҭÖ�'�?:��͜��{T�( &�^,3\[�v����|�������:ϋ�k���Kol�,��Ov�����+8w������gW��0o�!�lهW�/�)vo5�m"$���Fh�H)>(E���;�R�]��Zl�6��у�2�b���tX�mfE�?��\M�SSO24�M�=�Sƴ�?<�E2-�I�KW����B��u����k�Ga�>�M��(�N�Ƕ��;G�,m^G
ؑk��y�	��IU!tK�d�W���Y�#(n�P��'�rH0��\0{5,`����}��[q:@-��Ǭة��e� ؓM��k��%�>�kn�-�dV�C���C����yJM0��.��z�2�qŔBO���K��J%4Giҙ���J S�
�CB٪�SMp�������I��4�'�HA��!$z/=]�0(���vUb#��Mexu2��u��I8$Q�GA&���C�`D�UBr�S2�9��.������E�8tuu	�N�8��:�QǨYweg�J���M�K�@|{ڟ�?e�怓�����|!��+����,ץ�TW�ak�5���݃�!�c���������^SL�s+�ȌI�V%�I�d�]�&�3�.�qR(	���F��y}H	]w�;)h���i}MuU��.�1�R_&j%
9b�q�0
i$|j`��L�ȡ4��1����l�⌶@�i}и��S��E�7��7yh�8̳\���ED��1���qva��WV� �������������a�����p�Yъ�#��٥ȅl�@X:/vH�x�l ��@O'&c�"n�=s�2��ΰ^ZDI�ћCU����䗏��^�4u�f~��0~��X���LJ<UFR��zB��ȏ��K�/-G!ǋ�:e^k���hQb��T��gޑ^ ,�W�@�������5Y�q�`-�|-�h��qr:��(*WG�H�i[yW������=�m3vXj9��@���~eREm3�Q�����6hIJ��U�`#3ze'�'���nG�Q-A7��  $wq��{-@���u�GW�q��Y���	��ސ�/O�:O"����rin��~�u����R��%z�'�R�m���ܷݰF_��B��@aY�mH^��B�42Ҕ4�*�G�Թy'*�&�>�W�Z��6�,E��ꑿ����g�ԉ���Z41$��-72.|j2���q6�����]@y�<�s����q�-��j`*O ����	'��M
h�ɳ#Ph��s��5_���:�o�R1tyu���8�;��7IC8)%L�B�[Q��E�#�ԮV��l�5w�mv�.K�'�ݓ��|<�z3���{���z}�'�kEod ��L�F���df���~{5z�b���Y��B�RI��N&���j��)[8�?�&I������B��.Iϊ��Vh�W^�^>�-xHm�� �L��_���Ys9�P���"�Z�3�����#�T��07���}w�ѿ�����:���|�$�����I�b�-����t
�o�x�l�T�o��&3Jx�&�%���F�Ul� ��S��}�7��&+����[�8P�16��2!�x�H���|�W��rЈT��}R"��b�-�S�R��ё��2���@�U$�ZzD2ӫ���a�=@Q�G�,4s�o7�O ��_3�/*Dq���8��5ei��A+~���TQlD������i�[B�Ni�Ӫ`�M�6��0�S~�o��/_3�ZΦһ����*|��-�/�<##��_�q�Z��9g�?f�e���1�-����m|&q0��p���nl8�lGhx�r��}6T�����km�y���8 Q.yGD�����j}��{��R�j�~.����$�z:XfA:x$q<p&#�ʧ�ů�U���,�#m�K�o���ZS� ^��;�ܸ�ؖ���V��h��|�����+�u�_m�8y�f"Vx­���N/�|^?�й`�&�N��l}�ko�iٝ$�Q��������!&��r8��/i��3!�ƭ�y�+����L�9�%6��lL����T�䂞��~��m6��m��l�/������[?�b#��i�߹���Xg����s�D� �w��&�ɾ��g6#ߨ�I�a�6L�5��՚���: �E��E)�-i������� ��i0	x1��U��|b�A�?7`�2�	̆�[�X_a��.�mOM��K�s�\ۚ�^�X�<��q��m�h*�Ŏ<v*�D��Y&���Q3H�
��k�©�A��xQȟ��z��n����z��+}�$Z+_F4�R�V��^���^!4��a��)RYM,��� n�����.���С�ʶO�=��r����Z��QG����Ӿ������b1�#Vxt���4^p6|�������	���*��ב�M��h�B���q;f��``O�~*G�ՙ��Czw�pY_H���ϛoH�JF����h��(i�)��D���H҆nl��#��<:�N����}f��O;�:�5f@0�P�P7�gL�L��p����k�gb֔�"C�9��$��9�ڤ��h���]��ை,�j��%�3NKS��⚁1��ᰞZԥ��{U��*9�/m�Ƿ�g�##\�1�i��E_�o�)�q�۹�tk�UT2XMԯW��^r�yT���(J"�et���:�A��fE�_�󻒾.ſ�=��^_3Fy�%TN,�q2��b��z�$�1XV�7��8a�fx����f٣KDU'D�0��L{d�����^M�1��t�����+0cFL��6��Gj$�KK�����[��>��q��.�.�'H��i&L~40�x|�l+�v�2̸���{��&�es�ʋ%�������c����-�m�D����r��\�-��W�e&5Lc��O~v���"��q��x�3��benFl1#��m���ÂJ��@�����߹�S:P���>�A��j6�{Q�����X�#Y���iG�2�@�j�C��l[`� ��F�����ji�S�d$��"�7.fmm��t�Ox�-���^V+��Y}���8�2msWwD遲�	n��J0y�<iu���-�5���+�M-������A�%�Vo�?4S��9E��_=��2:�����t�����$3L�Pfal�����RW���S� ��`}�6@��$����VI����~̉2��B�v(b�l1�o������� �Zf-��J�Б���E�׹��z�gO��"p���_��w8�F����z�zZ|Ow"�,�!�X��G��T��4&Z�4dޣ�]����������0�Rc�yƦ��Gԛ�Њ5ć��ں��L%f|ґ�M��exh!j�x}a�Yc]3W5��a|�*��9�bh�_��f��F�ӽ�D�Z���:�E	�l;(�Z_��{�
�R~��������k8�|Я���<#C�O����s~Jr �4{o���^����b~ϱ��_'�ےң�|ì"�G�w��%s�:#����D4����2EVg���'��#��WI��|��ۜ�Ό@�*���lpo ��3"Gbn*b��a�͒e:)��J���e�'�+�Ѻ�2�9Q�|Ɖg����cf�ڒ��n�
�:��hd�٦E�<J�RCq-��A�փE
:��Ӯ��2f�@�8�aEVA96m��r���诡���M�$���-eW�_��+�I?�!!�i��O�'� ca��}�	m�.f�v�LA�T1U�%jr:M��u{�g1������v�=�g'El�	<9k@=���?�F��]�B���u�^�Z�7�wC����ɿ�-$�Y�7j9�������K�(�j5����^�ε�i�?�P}��S��Ca��X���,��(�����9�h����,F��K���2\�����r���K�n�G�8���-^Z���$*
#�����Z5I'q�ށ>��!�|8��vqZa��3�h#1�!G04OŊ��grl����˄�|v�c����PG�9zT F�Λ����-
$Du����}����p�kpo���<9�	�h!
��u�WB?&��D�$I���Þl��fߙ'Z��|�Yp��Fx)l���v��.�,\�"{yJ���f*�\�����o޵��#���]~O�h�ںCp
�n�b�G���q��B��*�iHK*�ܴ!�|-��&���^�ŒL��<�s��B]���Y�:��{��xa�}�E0�ڝ��I�V)���h�HQ8���'D�y_^q�خ�z�55�-�|�`����z���k��i�v�����C�e��e+��d���Zl)7|ˢQ����Ǝ��D��-�2β�p��<�K�/��8[�_�:�"#.'��Rڞ�:���D2�מ���J|w�J��*�������ڃ#o�T�ѻ�B�C)������`���O�N�A+�zjz*\�iI3Ij(�+��2���S��*N�����&�b�%6��$m��4��Ò�e�~������K����J�n��s����FT/�-D'�Zb��͑��K�H%^Q��g����^��l%��R�_1�U������k�,�
,gT�B�
��ڮ�bHd��B��]��,%������p����3 �ֵr:	?�2����J	N�]�C&1���&����ơ���4�o°�ng/�P^�+��B���Qa|����TN�Z���������|��A�-�D%rd��x̽w�i7�B���]45\#kyo��	9�[~J���UELj����~_�۸���΀'{W˔�)5X��1�܀q�?��k�$����(C؞;OQ�\XQ;�UR��[YCJ���������LN���3,����i
�n
I*WL��p���c��2aEsd@���׽J�ð�P�����~ ������a�(��def�Ԓ�AVS����$@_ww'�u�D�z{��`AҞA<���y���mŷ���G�=��a.�����O��:�_�9�!�2V}�+�k�c9HB�t��Ze{Gdi�z&�B��D@slwu9x��k�����uj�s��}8�9�Cg�u,�;O�yJ�����?�ζ�N�`�12b��iD�Y��y6�T�D1�>��Bg�%��v�������uVb� 
��c�㕾6��d79��q��M��8�۵�W��^$:�5�{�,�	E�</���I"Pk�Ų��4*�c?�N��b �wD"��j{,MU�r�9�z�ȫ��c���ٙ�6j�WD;wW^�����9�-T�2K�4z��Dϳ�������B�;�:�+��,�j�ڼ�Y�ox����ǔ�mu�p��`�@������u(��Ӌ]�C=�LR�Z�ް����L8����z���M1������!o�]��Y�&	�HrH�"36�n�������
ށ���9,�(��?�g"�s�v+�E��aJ$���Ö۽������}�'t�L�<T�ғ!������E�	` ��7u!z�\ɜ���`��S�Ъ�d���� �EӉ��NȘ|�_M�L�D�U���"�	�/:^Ǆ�0N�;�=�<h��� ��ZQ$�zSƙk�XOZ�G��xE8�2��ɠ▟�f�WJ����w�k�~X����3�m�$����ac�98VkS��������$��xTM6G�	$q��y�[���itČ,��wl�a8�f����H�`���Mn��Y�}���K��>����1�@�>�ң��������ąY	��k�Iפu���o!�̎�e]Y��H��D �������������4�s<)��樲���7' `��=����U�dO�͏H�o�����I�#P��-{#^}�M�v�t̡���ܱ(����d��R����y.�F9l�}�?%�/HG/�̯8�G�w�M�O���:�)=��X2�-�����A[HI�w���~�����F��ʎE�K\ߐ@�-�������8��	��z;�=K}��7T�:��j�yz��nb�n�H�{F���2h}J)E���/����4���{ܯ 鬒�Pj��z���ۥe���U�/�,R�,kH��X:{R�:l�JAۚ��8&��{�y�]�p5|�K��Pw��[�{u�1A��J
^�M3P�@)C�EI«W�q�����85�54�Rq 	y��n�J��*���-:�:S~�l6�������OQ�ْ�,lb��@�{��F-�\�	nͩo$�'D,xdKR.�J�
Ri��`tOh�&	�)@<
�X�uFeQ�sʆ#��(�/Ⱦ���\`$z�yI�U�l�^���A9�a|8���l:%��@&�/v�"C[p��,�[�����?-.�ӫe�:��n#�rO��0:��rH&,m��Q�����д>,�#S�6{�~Y<K���UX&��C~W=C����c����� �IBc�<u,kg��᫁�*�xX'+A_,M���A��ș��9IW�ȼ( ��m�.���(u!.�u��������i�>W*D���B¬u�0� g�ߠ��t
Eߨ��ҫ&L�=�������ë�q$���gN����2u�cCC P�l������♡��P���a��Һ�����j��)}v�ɍ�l�g��5K���T�I=GC��yL�|@�0g<?;+?�?�p�~�O��������هX�gT�)��	+��G�YP�ւ�aVX���2��`���'�}�=(��_�T]�a3M��w6/tkw#��`=v�7��ͨ�K����m�t'�ו8�>��ꮎ/����f��D2C�ΌM1���\�׆�S8D��P7!���'<����$ܸ�ק4�-7nu����S(�`��.Fd�����k�s��)�[��|ಈ�@��3���Iۖ�3,wP)�er��l��Sh���V��N�eKU$EӋ�;��ŀU��<���U�1x�w�Fgz��%�vmSQ���iY~��uIٌ�`���L�ٌ� SQB��2�����F�T���p�������2�~�W&eI�+^��inh)�:�E�AV�}h�63r�p�zf�q:�q�#'��6RCH�(0��#��Á	�d�oz��-�E�w�ȸ\�ȡZ5�c��w�dU��|�I�5v��\�v�� � �-D�E,=cC�i���6��'2Qq>L j&$K�:w3lٹ^��gO�u��KD��'��(5QKWē�*�?��}Si��@ϟ�Ŏ��O�d��2�b�$�w{O��8Z'ǥ<x1#��&Or��\�xă,��6F��38�^��J���C��ݒ5k��(^����Pi��� ˒.�h	9�~��k���M�5G�1�0���C>j�*A�a�WZީ�'�О����u�R;Se��5�~^;2��%�-{��e�.]�|8��`8��xr3�[?M� ^֘��uy�k�#-�T�a|ɗH�Y;$�3�(uvҏ�\���-K�~��͟�0\ ;9� ��*3��;��k�����pi�7�˟����N�F9��U����5���|�7��$s}_\s)�&�l�sm^;#{X༐�U�St��i��NMA}r�|��^s�r-햬���I��a�x^�GY��ђP{���=�����Y���^+�]Ϩ9YO�n8�رA6���1�l�p]�����D*J���9|4��D�h���9c��rW9��Y�ִ�L�������*.f�Y�-�X��X��_��{��ug�N�h�X�ȃ�׏�+�����R�s����2UQ��y2b��Xm�D��+�,sJ����!
�m��I�n8��s%,%E@�c����"�e�D`X@��
P<�X�����~�j(9�������n@� �ε�`�&U��*uߜ��G��=ү�#у����6+�f�}��?�{|���is�!2)IU��&�es�H�&6�˱o����fL6m���T�?#��dS���=V�@N�&>@8�`%��~2-w��w��#��|,Q��0�{�x�O��\#f���A��C��˭XdP�Vd.�V���=�
^��%�QQ�%��$�2������w�+�r��.ِ��e�j?�Rh8���`�{]��1�D�bbڜ�z���/2!�N�J�g�7��/��D�B�Ee�Gm�W�j��N�VNI��Z�!��� f
#v��\��Q����o6N@�Z�U��3wT�"� ��ND\>Q���k 6)-�/��j��Za'��tQA�H�_5��h'}�K d�亠��x
H�� ��]C��3�٪�XC�����'�c����|=�^�m���7�S�&�^o��(�d��_n�P���>>�,ș�4P>M��V���E��ν��k���M^�����T<�e�A�2w}�3��i��C�-,e����ԟ$��Z �cA~V0R]�^��LS��r
����V
�l��{tV��hS^`��u��'�	��0�<��<s`S�2w��륎7�"���8�i�Q�)$��m�f��E{�hc�]3�G3}��8
iy�����Ӻ�N�����|��)�.������S29���w���䑥��p� 9}b$���Ț�$�{�.|��=����]�����]�h�1K��cnџ۞��z�J�3�0tr��F�*h$� s��;=-�YRY䔧�8�����:D� a��SG<k�MfT��|�%�^C��!H�öv9M��s]��^G�� �ڛ��X�(��V��V�C�ǟɻ�����w��ZMe]��Xd ��h�a�!!�<6��S��6�;Nt��2J ���t�����D�)t���#K�8Ys&V-e��.��X=�E��u��\,O:�\!��t�s��CjW��u�h8J�D�-�K�dt'�"�QaR�w�Ϟ�aމ�:��]�M�N_��/��*#f%��g�A����O}��'�E�T3����a}8jQ��:vsS���E8�������L&��C�k-'��,J�p��1`�?��dk�m������%kh�Fq�6� �Wr1�+(A�!5�:��g?����ϖ��n%�/`�w�L���a�J���l�� `�&��)�:��&{f?Oj!�;:{�%4_=0�s��o�4) �+Ǣ4I�����W�CI.�L�M�*
���d�Y����j�w�ë@����A]ڍr���I���.��
�q\2�5ʤ.{�Wg��D������c����{����%�QM�'/8�^�~��T/�")�����>�zg[�OݣФ{�b�m��I�v�I�Y�.G�3=`.sث���V�l���IV�����~�!0��gQ��O�p�*���Y}��&�'��.q��&��y#�<|�y��.��i��(��{<8��w��<WF�-{�NP�����P�(�R%��ub��;�C�2�К�����cg����'X��7w�(��`4�l,�e� Bֺ��#��j�L������ӕ����qY����e����b��6�n ���#�kn���2lZK���,j2zQ"�u�ˮ+rT�)31M�_,ruSN0W���E�U���L�[EȷFɰɁ�y!�(��&��DD��Q�*l�k�WU�匢� 6�x�o��4��9����Dc.�&'���T�U���g��i�u����~�$�ȏy5���G�2Ϋ%�3C�m�!<߭/��z���f
��4��|�@�L=�M꬏&�v�X�%�c�^��$/�7{}��9YO�:aF������{�@x�s-��A��q����b��9��~��;�%�����N��Y�P�P�ڴ��e0x+�n�eЉ�h��;ǌe��ٺ�K�VO�ĺ�Љ�ޢ^Ōy�<�Z�������Q��˻�^$���N�6�J��s]
�$�e�^�Ђ����!\0�a ���m���[�����8�q�Rn��|��s�/0��͕`KS߃�$f.�8˹ۜpM)����P;7HUfHXcL�J3�8��1� fB�r�R:	�d޲��	'f�r�o,j/����R������gkC�f�V	A"�g�kC6_���Y�����	zr��s��e��떞VA�޲:���r�}j�/��w� A��a�L�MU*� +}�Q����ܯߺp
�S�}ep�5?b\�V���O��~�p�0$4��0]��zz�yo7s�b:Z�dRAV4�ìl�Yx����x�0f�5���'Ʊ���h�J�������<�'�u*��[g@
��O??�&A��k$h�[�~��j�9�W�p��'h���O�i(#^��-"�!�''~�TΝ�� �÷�����*�]I��TC�����s�������5��R*�ލ9�����Sߪ�n�
0Q^,���5����5My��tF5`ЍAnB�ex�%��Z�����#�$���E���b{�G��Wpf�n]��`��/G���ށ��Zaﺟk�g�g�e�����d�[f��fM�e�'Y���������5�s��)T�� p���V�v,��
@�I,�n�hv��e�q��������=>Ӓ ��K��Dt�镣�y,T9<4.̯X�Hb�)��E|��ǄlRee`=�	xӁ��]< ��l싯){d�rT�by��?$��W�΀��1�䝻]��n����3�����=�������� �S�����?�B��Wg��@f}���{�{"�}��rV	����w���PŹ/ok� X �f���s��B���#��	�R�8=�_b �uSRn�I��L�j��t���]Ճ+��3�G����v�ung`�Z� �
�C�gO��­�`�
�/��I�+��,�P���l��,S�~��	�Ɏj"w�0i_W�Ej��� �b�3߈�gq��l����Zb`� 5����4i�8�S�r?���X�ڀ���k��͍���=,�/j}3��J#hi}|����ޟ>��p��/^�&cdA`y���1�y�I^&�v��U�]<y��4�F��5�ͷ� ������N��A�"��]�R �;� yX?��'����*�9O�4��&?bi4m�&�YK3B��N21�/�a�3��Yd�2��:k�}>npc2]��H��4���`��!�.Z����V�oޅvM�����V�{B�����k���gتGt?��Ш�� '���Jߡ!�eEu*��;Xz�j[�V��r�X�Q�KE������ E��I��?�����K�� E.E�I�����V,斘�PX�A�|E�l�y�=:=`�"��~��l;�ɀ !�=�m?���w)�9m���=GPG�7��"�g�=�£���ٙYS���8%��(Q��l��� ��w�N�[��T ��x��O(��˭%��M̤�a0�a�|��G�������2��*F���mVp�\���;T"i>��D Wʘ�4O�h<E;��r0۾�O�a�����_q�(��a@|c`8�^����Bk��m�+;�^�f�5��5��#��}�����Kl���Nם�"4�X �p�]R�u�D`�����װ�2g$^�}x�!����{x��"<��ƃ���&$W�1���֑��P?*��o�8+ Ao�xÇR�ΜP�O�&ϱ����E���uW�"m�}�/��D̗h�Tyl���^5!���;A{�y���We#W��X�av�l�ˮ�Z<5�V΂��>k�װ����A�5@d;hS��o �~�!d*�R�F*ͭR$s_d>weCR<��!�g�2�K�}���ż����BX��uQ��q\Ur���'_.���MR!�,fa�C���5��Tm�JO<M�[z~�*�Ѩ3�8O;�$U�B�4&�)�#�t�NC*��Q^�b��Oeꁵݓ�#�G�5?�:V�m�/��3v�t;�txp\��9+}��CP�NOc�~);`=G¹kzh�RsM��LTe}��v�g7�C�2�ʲ���D���,"��Jԏ�T�̄O�w�ܱ5�8Ỿb����Ѥ�2����Κ$�!�7����
\Ջ�9��'ʍt��$���;3Ped��M>�3�(L�d(_����e���4CMɋ�{^�>GwN���:Gp�J�F���Ж����T��:Z�7#�Y��kS����m��f�M���%uD��	�O~|@��U[�?�>�4���"�Qq���s=P�ɦ�#3R^��&�#��-��I2���i�3�ܶ(?�tG�&g�̐�G�RΡH�2�5:B�H\�-=?���Q�+��R�ŎԵ��ä��?Ev'�*w����I���c� 7�L_y�M�%<^�R<�o�O����r��� �}q�#/C��o�ft�I}�3�ᝫU��t1P�gc8m��Y�M#!�pPMx�0�Y�x!p,O��E�|Y���5`���"��8 !M,��J��5�����ހ��e3�Ǚݒ��#�O�GI��[<��A_ĩ�s)���C]�Ǣg�Ƴc��VD|�MQ�%!ss��]g�����I�g��4�����N����8�>��oV�/a��I �e=��q�v4uB�WEƾ��~�9%Eh�L�*H��B���K�n�n�ߝ�={Po;i܂���n��0�\�&aDD�vb�Q�JhG�'∰$}��v[^��i���X��d~��5�\ѯ�C�e�&��?d�V��#�ΡD9d���ː�鄍O���T{O&SdI�_�,�Tm��R =_�*xl��h�%A���T�ϐ��yd�W�;��e!�p��)'���w�1^j�Zoi�gR��޴?�Ӗ2&(��w�J�ɿ��Y!q�)���Bmߘ1�h�B��|z���+Ny��`H�`�JѪ�x��̌>�&3��.w�~�vWR"�[������"���[�����)��vW�d�9�A+�"ۺo�P�1�ZU~��O�t�n���4��;z�Ωq�K�~H@>8x�|�ѕ%�K��8��<
GM��%ebYfB�}:3<,��ۓ.�箨Z|���45���KfYS�+c���~I҃~���f_�A���G��2j>On�����D3F@��}�ؔ_%5�*:PzN��=A0Y����y6/:RO�^�f!U�o��;v��U��c?���V�z�C�P���K�Z�����&�� >��g���[E=2Z�L�ގ�"������PX����>��U���K�[~��S�t��rk�D$X��Ըf:T���� �1L��+ݛ�#7�e'��V���7m��!�X��98���ނ� �׍�`nE�?�=�37-�7n���	�TS�y����*�'�"�bH?8BH+�ذv-�>� &w�ި��}�ǧ�989p��S�ΰcbF�{�JT���f\�5���2��M��j����3��	j�T�K=�x��**3���T2\��i$W�6��ҽ��K�cJ�C-հ\���bxo���|
��μګ~ٸ�t�����x�ĭ���յG�t@���`a"!�6BL�s[���|�
�Ϲwŷ������qd�����Z��\��ȚL#�'�j갿o�T�s���F�U��(ô� ���#�pt��@������js�qg_lKT�[G��S�E�@\�YD09C����#�`����4��fY�2��������e5�d��X��j��np���I��	K�ڿ�>�C�����"����a�M�PE�[f�t6ۢ�c���;y�Zr�!��aL��������f�;�``�.cu'����_�['�2�c}-��;�o���%a��jw�/�=&��HeIũ|
V�!��f����2<���m�}cO�5���ަ=p�8��+G{��d��/,��}�J����{��p�L�|�8A����y".���rV�QA�a����D�|�G61�
�LR���A�(.�"��S�"\�M!l�V�ڶ*ʨ�.�1L�v_�'�OIC)��$FvpY����_��V�l�wR?��q���= �~!���fl�m�=P��4���`v0��p@ėk�B�!3�o>6imm�״�X�m� :�g��|Ց���t��DՃ@Yc�ָ��x6������������`�߮:�sjrn8��w�g��=��{��el&5���I�3��;{@c��Ф`��(c<4�KHygY� 3��~|$st
�B��r�D~>f��!ib,���qK�G�H	g*�7@���Hÿݘ}⿺a���y`�D�i�i �liN��M��s�S�b����Jɦm�k��:>_��U��_/��1%p�K �:V�Fq� ZG����X6	�u�2g��0�׹eN��y���N&,&�ܦ ��\9�����2��l>�3C�������K�Δ�c��v����(>߉&�W[<���1��?��^K�����t�����������O�R�.1�d��ؐ ��O�\#�q���+��Wu	�Ɖ}uuN���r��c-{�*�qڜ%���ޣ����Ժ�(#H�W�>˛��_k[/����z�j��>>�G��#P1X`�N�e@��F���)\�;Bb�nﲉ���k3��LP"�����V2n�5ʹs8��⋑����G٤ނ7�c�4�''�Û����g#5������Ǖ�yqPe�vqkm���K.�L&K�C���_��*�5̮��ύO�B�X96��
Ԩ� N`��U$E�����.��8bz@����ɂi��X�x�� Pޡ�2F�uV����#e���u%����Q�Xm�K[��0&{�����<�'�g�od���u4oB������\Ð�W�Jh�K/Q�b�غg�'.&C"����$gc�$F
I��U�,��n���r&�g�mV0A�Y�w�̾p��[B�H����۸e�q ���柙N��ꅷ�ȏr}�G޿9OCZ`z�2r�B���N���\��E��y2��z�5B��DW�Tt�9qzX ��6��~_�b�������Va"������N�|���׀T�2�1o8դ"�	�GL��#��^�F`�"MԠ�W�!��05&`[Oѧˎ��*s��N�m�H�pa{��;b	�v"��ze�=�pn�j�v�U0/���P��G�e��l��p�&��jK���h�<d��5�:��N�7f#�/4�?����4ZeL\4.]An{��SW_
��/���Dx8 ��p���,޶;n�}��lI���#�����9��Y�����̘Iʩ���pSD��,������b��ne��������:��%�ᐬ���^�4BW�g�Y
�M����X�x��02@�9V�q���i���'�@d���M�;3K�,��up��u*kɺ���ej.�t�oP�9��J�R�����Ut)����s�/X҄x�AC�w9�4�rc�������_2���tφ��;�K/_���Zj~0���,��5����)���Z�HBr��hW��ܨ=��-�%� �{�S7�A�W�'���u�8�p�0��Y�a7zS���������[I�4u�&p�ԖC�QJ���%�l �/sY-~�q�U����$\B��n��������6�:>�a0�C\|uY����?ǻu�&i��6��n�|QY��x���޻����yc#�HәC=��m.{�^h)l�K����v0�&����yv�Շ�)�,�QL�J��MC�"偏��zw\����#�ऻ�%�V۲
jo';.�T�d 	���7���X���+�Q_>B�aJ-9@�r_� 5q��E��~ߖ����uW�D|?϶�6�b��6���=Ke���E�<��7�ʕ�R�������@Il=�|)#�.{���6��Mi���G�R�n���&��p�����čp�$t4��N-��A��y���S���������K��";�M�9��������o�C��� �����)�@0EX�܀1M~���ꇗ~�ǅr����+�UI��O��#2�Ϝ�)�#����LcR�:��7JH�uҍe7 .����S�&/�P�꾰^i��F�������\0�u�V<�\���w��̜�4�j�� 
���+3�nP�)�ݫO��ʃϘ6�>p�㰧u��vI�K�G��+����{,֚)�t���fE����=A(��2���[�̭����3�=�m����t�����k�(�.k1��[x��p�4�m�{���xMƑ.IGFSƂ ���铧N_f�t�%�1�����s���Al���lE��r-F��c��C�jiX�J�
����>�˶I�	Ff��Ω�@Q]�y~'�����?_���x��X�3��Q_mU�3;Ht������m�@����v�4��NO�{�~G�`k���,��v5��Q
�5z ��љ���6�؀���i2mo}~��z�!�>t0e)���7�(�����E��ԇ)c�5B+hCf��/�~k=�T�t{"��BǃGc�a@w1X���B&b����}����P��4$�<��L[~Bz���+���L\mҙmi�ӨУ&�_2���=�-8������t�F`��;�#��{�@s�d91�
H���hX�j@��p�'�)�I~�՟�[=��}���p��H�"+�gl�%�l[&�8$�A�u_�ڠ����*�V���!~�񶾞��c2��+��	}vp`�_H\���_
VW|T����6�j�[�f �k���Ut���'~��^mcͿT�A��Ɂ��@��0'��	;�֍�<��JP��G<���g-�s�]��7��XR?*k�Wė�M3�[-Ƿ|?����Rb�v��o���3H�k�p���4&h��R���b�gT��^gSR�����V6����7E�!��wc̐�h��A����R�� Ң�7SJ���e�Ո>��A{��b��k��h1cl�hF��:� -�F��{fɝ[L�v���Q�/�b�j��m�����;K������bSc3H��lf���3�$���ɷ��O]�!L�(8����Vs̠��AK���)�o��h��ꪉe=������qˆr\���+]�-L���`��ԃ�O� n40���h��Y�6�O��W.`9^���.�+�䄿蘬 �M-��*������9�ag	V�Z�8��w��S����]ԁ���EN�����1��m.��j��f����Gd̃����H�JOz~��[ʩ�J� c�#
� z;�[>�r�d���qױ〮�ت�wA��z l&���04vBd*R�������6�|Y��8�S*�q� i�ɚ��97J�8�W�WD�>}@��j�8K�(�����x4|�/���NE�6���ݢ@����
Q7h=���.��yTv([·���t���?6DY6'

�jIG#Ԓ��g@ sYy	}��"p/���y��1��n3��@p�EQL��l��MSg�:��\R��&T4�U2k��Ҿ=�V�f�gk�A�[ �;*/�-p�U�?�Aw�
��s�YU�������v\A�I�d�4}\�1���u�7���?S	��^I3hۨ/2�1�C$%ۥܟ���j���䕁��=�S3o�BMi���T&P4��5��x^5��u��i԰c��<!u�=��"e�:���1�b5�ݝ��
ۭ�X{A�[Lɗ�U�p�:Y9hF3=�Z2n��FZ�e�o�xF��Һ�����x���NȬ��_1���l�p9���(��|�x�����K\X�,S�3��3�b��(��2A���L+��i%M	�/�ܬ<�oJ~����K-bO݅�r��{�8V��>y��K��ʐ�[C�p���\Ts�� ��H�`��Ґ5���r=s���Pa���J�
�9�脘~	۟�=�-|>�h7��Ҳ�[�HOˮ���9�
��6ю�Ӱ;[d�Q�!�UDV��j7��V��R:P�8i(m:���C���旽�Q%��ۢ٪��h�V�g�N�$LH���`6Q��h�_�uS`*��ȑ�+aZ
,�)��j��v��3�	�����p���X]R��Cxb[9�rg�Ca-C�K��H�屩�P�y��30��0f^H.���x#;u��vzf�j��,�&�����3Q�B$].Yzpρs���"�M��4�x�\=`��a���]��5����]/e���D��)*�d�~nZPݖ�By�΍��K|���kg���Q;���}Am��j���ӎ��Wfc!�D�ڞ�Cd	�K�kT�>]�GwRR�(����^fW�<~���hl�V�d���5��*�E/j���d�����p����1ŦW+�"�r�#.Mb��Tp�쬀kc�S�Uzbp�F=�G0w�ls:#�8��K���a3}��+��U�a�n�L&�VAgB��_*k2l�S$��>�k�h"�<
%�W9�z�C;u��g��?"�>ܖ,���R5��h�H��: �p�Z�AjLN�����Յ�^=��H%�Q��f�U���_f����7�n+���}���3�����9�4A�yC[?Y��W H*�Y>,>yJ���Hxw�s�{l+ �s%x*Ջ�c�]�q������ZeH����pe����B��%4�*H�7�����J�� �Ԋ ]D�g{P����gJj	�|%�6Q`�!�]b�|�ΐF>ca �!����z��Q2��e,0o��/���A|}z%}�@�[xy}Q_2��J��§��P����Q���\qop�7E�+�j��_���FMA�H�D���xrԐ��4'Q���d�ZtEω��ݙc�h+��0+�T�Sz7��W�:��V3	��R�������_K�9��L����4�^����mӔ�hk���Jvզޠ�Qn�5�&�[WZ _��8�y`	�.��gh󏇫JS�� ���Cx	��G��� /��_�$�7����1?y 7D �Dsy�W�A7k(%��qu�J���i9��y5�w�@(/�{Q�Bg@p��/��|����?��E�]�l^�ڇW�/���FV��(rhi|r�7�s��t�Z�f ��",����J�FN�`R��^ܿ���y`��c�`U�I&��������������0yi+��{4��jIY���^�E� a���ʘL	�fP�f�p@�ΐ�E���E��Ojk,�J�!q}#����?�e�h@��*MM{K�^��|N��X���
�V�[T��t}Qb�m>�qƁ[����eM����M	"�JHS�K7��5X>��2�x�{ �~�c���Ro��]M�P��L-:�qF�v_��"5[�>������~���v�'l�zb��R��E+·�K��<�`gZG�3cI]T��uG��&�zY%=Ҡ��r�#<�:����d�5"�U��>0��r-;��6+.�������@ge�c#�fЂT'g��9h[!m
в�&@��ڰ�|���s;ֽ��~�����e�Y��,I�����:�kg4��s*��nO�x���)ݟ"[r$��5NXjٯ�n��k��" ��dX��]��_�0�l�`[�*��.|���E��\�{̈,�M6���eZXm��y���?�;8��A�san�*zO�I�ۊ6bP��qʜ����Ë�A!� �0y�&��ٸւF�ʐ���f�4����8�,�_ui�#R��I�p2��~ATN�\S�p��X�<�	���;W��vz��ݕ+����{���1�v�1���;	Ϙ���s��<����47�ÀT��φ]4|�!F_S��I�c���K�(,��$�R�Y�����#�0��})�VU;���a4o�7Y$:1,�.kwZeދ��`Jxm�)�����(��"���y��Bi�d�~Q.Y���6汨�*�gF�`+Y������'W���h��v��:���i~�B�4@B\��$�G�.�ǙH �]���~�OQ���=e:;���G��c�9ϸ��me99�PS�&�}�%>�
R��\�E���|6��)fT~e�s&:��m ok.�y�t/ف����3W���%!��v��RU$r��L�1Ik�RqR7<R_)�1��� �q�́3�Ğ����t�j�)Gٶ�2K�wQM�l�B���~[@�'
)���ù6��O4{��l��Cl��l�~�h�Ɋ$K��|�~����Q�H����v�)y�J�g�UӧH�z���48䧺�)/�"�^j��*��悜	H$�&a��ٯ����[r�1<�W��:�3�'QȆ�a��Vȷ�ShJ�6{��vH�Z����!<�x�VR���"]��%�{
�_�7P�sc��%���}γ�,��ד�9�em<��l�E+�.آ�/�)��(����>��J-K�*���\��|�N/y�*�}��� ��Q �?��zY4v��'d�}h-\
��A��$�>m����WAș��vY$T��3V��$}LůJ�dRЫs�����U.�p�u�|�'�|�|Ĳn���i~_&��^�,Eq~�,�{�%�ux;O�q��B3�Of�1ƺ���m�� g��n������	6	�~~��y� 
���ַ���gb)���O�+���l�l_r,Bb�w�t=�E��*$=]Wm+5���}e�`&7c.g�w�w�&C:�hu�e]ۂj��^��pǲt.���e��������{��
����#ڞ�^�q�T�����č�H����f�-G��rg��f�S��E�n�#�;�I����3N��p4�K;�J�d�$6�*K�s0hݓjjΟ~�����,�{�L����)F�]*�d��Ը6���1~�)�]5^x�`�~i��ݸ�0V��8YO�D9ij����NGt���QX�0|��8�hW*��Cͨ������r���\��W-,�����OVd���3&C�Lt��O%��N�I9����o^i���r�pז�,ܚ4A��4!�l�$�4ER�JCk5xԷ?�W���n�����N(�<��6��γI�x���M��ך�Q>M��z��\Z>��W["��G�c�KR��eK�A��fy�me�C�����g1Y����C�s�7U_`c	ʒ)��p��02[���F��yQ��2#�!m��L�g�3��j8#���u	j\���bB��Z�34���6�^L�ڒ-��jwn�����D-����qɞ
X���J�����J���NEOl4�����mKS~�5����I
I{w��c�3�[���vD#_})��Ɣ���t�к�?���a�ML�s���>-Z�G�;����ҕԒF�r�C�xY=!.�2�m�͈�����W�(��/�էǠ�1�
�J���J��	�o(c���hW���}Rb��kDm_	r���4	��d��=�պOF��v]�oS���烂52�b7�(��:����ǲ���H�lC��q���7�t�ד�Ϧ_��)��]{�if=�3!�}��.�=u 0y�R��G�a)P��g�M�-��/�!��)=+����sN��`�I��#��A��c~0��=�_�a3�h�G�N,q���@��T�贎h���w�L�f��ev����Lb��U[&Z���O��[N�<�^��8��6%ޣ�sʵ�#3iG�5�)��DQ̱#�Q�S��(�ٔ�D60���Z6sR��� ,�ɠPU��~]:�:S�^r��c�v�8i���W�H��� Uk&߬5-G��P҂`@#뮦��W\�h���.4�u�^w���s��_/��dv�+U���][����O�T���e��ΰ}�����rx1ժxr/�u\g�Æ��0�i�E�y��`~�b	���W���)�v>It���g^H�I^��z?E�׫<��ˬdJ�B�ń#iZ�7yC�?�#���TZ�B~�O�z��ܽe�:%OS����7A��ǘ5V+�J�(�l�~� $8p����3!��s݅$�mֈsޕr�m�^z�7x)��~s~�,v����Nw�ڹ�8�t����/I��3�;���-AVb�Sqh^G��&$�ˊb�5��'+�_F��7���Fg�"��D�3u5^,�ʗDM�|z���]
��Hφ�@�D���lf��ɥ����KvԵ�֑����^�ϱ)��FLPQ#1so�%9z��s����{�Du7ꃉ�en"B��T���-�����֧	�����͡��� П�~��K���ѹx��>j�x�m�P�k�X;%<G����QR��k�U���r�a�j���ԣr�ʉ�(�PAx�Mc�����[����>�~��Q���هc�dQ'@���I��N�ҿ��
��T���D?C��m��ˊ �wI�X����k�V�fN�1����H-y�o�~M��iA[��}~ބ�������pi"��	cw@J}�(���57q(�o�f�m_��]Z��BƇ�:ݻ��육�����_ߢ���1pO�=���2�ʆÂ.9��P$�xhS��������Szޫ�Dj�=C�4G�K)G!7�Il,�Y�rv�j�M�& ),rO!�����N�A�m!�L��5��B]��Nր�W5�5ۓ#��o<D"9��cq�B7�!�����o�l�vr�ҡ<cP�������I!�(V��>d���:�r�Zg9޸$*W��VP��(��4X����9
��]�HS�/
c>A3FYǹ�@w~L��i�6ױ��V� }\gc`�u�\���"�K���Q"_6��2r�.�޶Lʨ�Իӣ��0��_8�����̕|S�|�ܥ������U꨷�����k�%��v4�Л� #ĉ��_G��,����m���y��e�����F��p"��]
��N0�Ѧ�����$`KF D�1n=8�y�j�"Ȩ���ua����b����ښM"��Q�� �x�2�x�%�;�&Z�cvcx�M��PN(�lY�~T&~^�|�-a�2`ׂ�j��Z3��^R|"��{OI	KV�(_Vc���i���?�N? d|�w�E�c��R�E� �Q[U%@�^�s�&����բ�(@T7�
��%�>�ч���uH�!45��g����ǒ	R"�/8�G?�`L���~ �+J�/��%�DqGU� %���W S�P�4�_&��po�Ǜ[w�9������W�U��f�l��?Wd�d���C�T&�T9Cz��cӸǥ���Jl�mP��m ��٣E?��WvFz�=��u�z`"1g|��������>�&g+Tհ��P���VS�C��)K�x�����M�`[9(����.��^���������D�}N.F�s%}~�`�^�̡fh���\�lWW�ׄ�\K��,iiB��6 fT�G�2��_�)N�&�PW�&r�S�}���4�\��@t}���UV��3���m�6��l]2*|�"K_wr�6�/&:̦�)�S�R���/(I�!��at&%H\��Ԩ���ob#�|c�(���d��ڮƂ��21����}��R����{�����7m�,��qB��ۮ'*x��<[`��#�/Ր����NW��A��1A� ;��\
Ӱ�W'w{�����t��AF ��mW��0����9w3�_��~�!}����17�	C�^&�VS`�yrK�-����=_sA�PLh���S��ˇ�����ؠI�c��4���P~R5������Y�s�� �׼��W5�_�L]�<Y8�TE���������Ps��Ak�M�����cf$j�.WS�T��}Q{>O��{Ot!> xVA�����5u�}iQy�M��0��5��=�0EE6E�]�o�˒}9呑����[h��UG��~ꔤ���(e�ǻB�.��^�ܖ�.*��L�q��gmu�Rڕ����D%^qE���J��G��@A=�o���o
"�n�e#?_�r���<u�x)�-���j�{G�
Z<�0�۹�b`붆�bзqOkh���1�W�u�:¸������&켼��T�2��OqO�3��qr�!�{��ӡW6vC��!p��%��;�L>��4�6Ǟ�:�ϟ3_����Ϙ��w��و��bl�!�>aRƈ����B��U��!\@�	%�1��]L,��26nh�ә�Hx��1jB���h���^���Rk��
���[����u%���f$n_$p�CJ�K6:]1>�R�Oe腃�;�ߓB���\k�zH	�jY�����|w��F��S��I��T� ]	�o�B`�]����[_�?���Xg>�k)�=�gw��(�D�Q� �GaU�DA������J��	ZѮ�+��D��h��ސ�4���U>�P�) ǯ>���<D[p�L���b�����Q���Y��C�wy⬐O`��V�y�`sm�<����i�u�,�mH��&�7u4Ob;�5��ܢ�Wl�<�R� �.�82u��0hg��I�6�@A{(Q�Ez({�&����ڣ)��}�X�2���~eI�,7ɘ#V0�w�,����W����}�k_en(HHxr���C�nЇ�L�v�f?�g0=z���P�C�x� �N��~�Vݢ�i�5�պ���?�����+�˥	|_NUq���K�]0�Y�x�c�/
�a�U鳿"/�=���I���+���=6(�����\������j16���sz+ʢОG.��bxG��NC�?H�-��,�O�~35N}>�Q:Z�(��?ӯن�[HP�����oc8|��%^��ޛ�-���J;�yk��@�3){)�e����/[,L��Ua��޽A #��h�>н�R��Q����-�Iz�pT��l�M���Ech� ���(֤�f+BXƹ#�H9��Ʊ㿾'�D�%z�å&����W -.�Iht8��ܻи��:.�B�{���
I�'��1����@��y�Kh���%:�&� k���)'Fȋ��@��jE���[��4�8^̂�"��q��sT<Y��g_v=H^�N����7�-f�̄	�^b+q
H����1e>Dn��C�e�ۅ�g�-d�59q`�\x�d�9���>j�.������Vk�ѵ_W��@0h[�߽֤������C5��O>A�Xq`w$V�����զ7L��5�yAi���L�5�ph����맱6TB�u�^>��&�	���$2-���k���R�=WT��2��ω�gq���l��6�Wn�C�=Hc�F�l�w����qL�}��Q��i)Ң�_�	;��C�Yq/���ˑn?����V�{��~�+���p�\wc?�ʲ�D��m���Tp*���&,H� [�'qJ*Q�a�zF��I�'�g��	�D{�����l������һ�^v���)�`�``�2wir��D��z>�C��	��j��*��P$g8�9���P���p��5�V�Y�M�q�̨���<�ܡ��u��|J���' 6��Җ��C��$R{���+�\4�]lp	�l����?���NϺ�-+B�g����� q�����_$��+�7��Q�D�K�<[�2=ts��E܎'>������z�в:�If]F�=�hڃ���H����j���ƚ
�<��t��1���[��^o��S������\��ᇎT+Z�'-��z�us�F6��{�p1�%7�ƍnrx�(^/�$A<S'b����\C,�ɥ=�Ŋ W����.�{�Zc诖li";[���?���ڊ6q)�'�lAm�K|�|~e����w�����O��Q
v&U�
�?��Mщ��܂�f�$G��,qe��C��I�c:29�ň��́�3A���m�c?f�v(4*�sؾ&tl�wʴ%��f˒���"6xֿ�?n��L��Ƌ���,K#+�SCv���b|i��84���E+�a���4���VT�'Y��*�+��?v��p���t�r����}��:�L{(�D��)UR��c�C#��I������x���v-{��E��I�~S���)�\W������Ʉ��7���L���ן��.�O�\���|+�⒀J�?������P.kW=`��dJ�#�sK]�vnh�5@+/p<���\�z!����;��6��R,��b*���k�&�C]�P �ۭ#���x�E@ğJ�|8��D���w:�źSb��g˭к����J�R�YS�yz'n�I��>i��^����DA��K��� R�z!l��Z����e���*|ߊ� �>�ҩ��ڮx��w¸�����qE�<�,T��-�\�R��$������~�=:�PKT����8�w7��p�9�e����Ų�ǩ|�L�c��֪��$H�)�c2����g鮼�l.�d����w��PYI��"����t��DՆO��C�A���L`��q������l�
5-]���f��@��J�&��09��!:��"鐊s_�WiX���LaX��x��W���F�LiD�
66�?�#u[mҥՃ'иtq�Eуnf���`y�#ȭ��>�>�lXA:���W��^3J���B�K,4$���<a�r�Ev(Q��	&�3%�$�V)$�_%�1}z��]Ȥ"xM�˵rd���]9(=�K��U9�l�MWA����z��f��2wĨ�ӉZ���=kU�=˦������r�/���ֶPy&���D�3Ԑ2U
�������4������K֍�]�R/�6�VA.?�ʜ�4x;:v͙��l�;1�(�~ؔcn���ƪ!��.�5��iq�Mݦ$��˛o���Hy�GH���Wk۴���J(���'��:����+�Ђ�U3�H���铮HL61����4��O �̌����uo�.��G�m�Faf0/�M{E�P�|+Gn�{XTʹ$-g�v~��5������~,|1��o֯�I�Nˣ���Ǔ��3�����(��(�Q6�r�[�y�����A�P8BV�ᡥ�&Fr��@���o-w=x�{!�vC>��.���	n���N�	���.�h�}�"7�m��>:��Cat�A�����U'؉wL�c���#���Ir��qa}K.To3EL��Z���!�'��t�J��ۇ�|�N��������r����(���Hn�4�`V�S�O���(�M�D�V
�O,iyg����F���bA�	�B��c�]�S(�5�.�O�����'��3����UK
�;ա��,D�~����`I�g��%�`zk��A<�ښL��2���ː������e��&4�#!`c?����aEY����~ź����~�.�|0SΞ��g�������B�R��F�C��5 ՛�������i���Y��� ��B.PzO�EPU�� �D�p����D����<&�Aa�r��}
�"t�%SȂ?`��߰j�A�n�"���W�h�글lc����9��bxj ��V����sX�>dʴ�L����ص�W�D,s�W$Z 0t���|G$������GM�=�Ƀ�&�����26�t��H�f0�\���n�Řf�݅�o���R�&�����|[�s� ��C��:���;��.K���^���r�F�4�Y*��~�N����ܛ}	�:J>�����-�ř��GǇw.���ߓW��i��w�z�d�]��n:h7��U�@;DMv8i�	R �"͍W�J*l~_��ū�u� �2�n.0���C�c�t���~�{B%���k|B�,��-Kn:���΀�s���lK3�����ao�>di�9D#=i����⣬G��4"l�6TTD�ON�la�b	�3�#!W`}�N���O���J�����Vw����K?�@���Xܿ�
�yO�E��i�NP�m<���$��y�>]"BH��Lt����dT������a����L��U�WZ�c�@�ࣜ�d�Q΁G��t0Б �Z�S�P(��Hmz,y[�9����m�����%2�w%�r��Q��e2�G �"��{��z+A��@���uD����rw��qj91݃6G+���I��䦃���C#��}jG%�z�%�u�`d,D��ڬ�߅=|/N#� W(��X�1�%Ih^4qĪn�W�!�̖��`�e�j!���O��C�C"4�D ���feô,]m� ��px���r��\>Zv�ˈ?���&�5}��k]Ÿ����͟+��fx�7%���bQtR�啍��ĞČ��r����h�Q�Dvd�}_
w(��H�H������x+�����VGa��Zy������p����SYV��.2s1�q._�#�^��6J�u���*�R��h�AQMG��\�<
7�sI㡯P��?�jW<��D:ކ�#�%��5�nS�!UqRm��� h3ߖ-?���ei��#.%MF[�z��@�T�A" 5=��,a.=�O�;��iVoXV�J"hx�@��xgtC"����ǉ�����e�V��}c��� l�f>��sL�n�
?�c�mb�����gB�%/I��wC%�$�\V��5]�ŵ_UL�w�k*���LN�j-�9h�}g��sY^ ��	s#Ԛ�t��l=�ǩ���k�j[6˝��0:�hp��vi;R���0�����_����B��7[O���{?duC1�������x^bgo����`��w�]�+<��*��^�
a#���B����]L3@l�;�0���Q��#	 켜���_p�MCi��[[��P�UJ-��z>o��c� _�iE���rJBA����ф���"�����y�p�?��~��bw�ul:0kQ�TL9����ƽ�7(��#�c '���T˵;�C��c_v�虗��Ɲ�N�g�X%a�|��5z(.�q�^�8�m�64eg�$�|6	��uqk�4$ƹ䢽j�
�Q1#�iL9Y�C8�)C�\�6�)��lTd�ab��AЛ6K�DmZ�3#l�<�e�s6��l�c^�UJ�(�\H�{Y��;�i83	�C=p=\����@{��{�?��q�s?z��*g���aW�Ʌ=�,�7G�'H�1�"�HsHJm�/["3�<�sj[�ٳdp����Ƽ���T�M�6GN{���)�C*��!ہ�Jl�κ�ɀ�7��� C�f��t���'�h"�]C_���$���c���?���ɾp@�vĔ|��&݃���g�s,n�(�u��U�>Q��M���ߌqKd�0dӶ�H��3ES��.e:�t�E��{����=�Y�&6�F̡��GA��Ο��z�[�͔��q�{Y���W�Q�6�Y����R�B�#N���7�ܞ���KW� ��({%JnF쥪6k��zy5%�x$+���:��g�x�ǹna���@���%�*`��,z�d�߱|.�,n��x�I�P�01 ���aU�֍#��$dX>OF��E��й	�i{�a'y��=L���� N����'v9�U�M.��f��u��H��}�z���!��q���5$ʿ�7&U��\j� �p 3�-��-U-�F��0Bn�L�8���A���9}�(�) � iv}���c5<�p�A��c��q��LH�o�îk����>���Ԋ�ʮ�҉A�*�<�b
����Td�\`��e�CZ��_j��ɬ��O��[��D��`�]�n�Z�P�N�{��Є]�F��x��e�6�4pp��dA⛄�4���{��f'��]˯�ሁ9_��|�D��-��\=3�B�|�e�T��(�Q'�� �5�r����1Vh���~객����)���!>3�'RG`�H����%R�W~��RE� f�I�ވC<�RZ?�~�W��*��H�t�;��u�Q�G���
�3c�	��?�-��}$'�M:�����0��۝PF��v�
�J�T��C�K�}Z�3z3������L���Dn�r�Y��D-L���Cݯ��ڟ�v��5=BH�v�ݬ�K����8ϜBh�~�"!����b�G,��R4��>�-�MT�!�n6���iQ<�b���:d�͕�����.t(���Y����!Ʉa7R�㌓��-�j���`�(;6H�rv	x=�4�X��y��<j8J����p1�'�4hVz�#�m.?0���b~1��L��\��.�K�6��BWҳ��vم���F���m`�F��p���"��A�M�h���< ��T$�t6�}��wQЌ�sD�М:�nH�����v�<q���;��?�@fZ�%#���֐P F��H�c7/�)ާ����޳y߰�W�O�<�O���ܰ�z�I�)ʻi�����P���1�4��E���2�$��_����m�~�&�?�*~�4�X0�a#+��Pt�otg��H��s��[ze-���yf+
�w�������G�t�h�ު���W$L�>܆T'�22�Y&�?A������&1�(�h�o�za��o���.-^tvKq����N]m�t��1�*�:9���j]Z���i�ֱ����{�@���F�҃�G�8Sr}�~��z����x�d���@���]}������O�;��D�� eb���b�(������M+n�[��ݺO�`9���Y�N�~��j9=d�[�Bt`��́���S�-��f��8BӒ�È!�_��X`�9�8���[�DYƺ�<����&A���6)	����J�ؽ��`����0��.Y6�����¾�ÍK8�4���LtP�Õ5j�k.����h��G�{����i��U�u i�P�S�fl�&lI0�ON�\��c��}�Сo���ڊ�g/�/�P�G�G�[����	�?]m�"�t��{�~��"����v�cU��@T���z��y� h�p￀ {�}�Q�L��e�@��u 6�
[sA�����mt�;���PX���&E���n���
����uA2���
���|u���p�c�����S�,>���һ��p�Xy/R�/�ƚ���䂇��J�#n�k㤄=���\�W��]���q�Fˉ��u�]%�ا� ��p���>�2���K����1�[��ֹ�q<P˷��yF�lj����;�'�4��OH�~K�TU�a��T��k�Wq�2���EZϺ�z��	��{3A���(�H��Y�V"F]}�<d���|h�."kzݾ�������P����c̓@0��||B�v�6�	$��~ӵ���pQ���j���(q?m��v��a0���0�����`�&}8G��͢�mVP�����5V�rf�'�a|�wĜ���/���u�j̪�W���.|�Vf?���	WJ!m��ʤ��Е���+%6���T��R`�O�yg�.1d!ѨI�Y��*9����]f?(ܵ�O�c[>E!(����f��jSk�r�`\��>#�|>u��I��(��Jb
ؕ��Vڈg�4I�!�iҮ��.�n�n#I"6�~�d��Y��}���Y'��h܀�6���q�nr�g�m���J�W��>���&R#���֐B(�ĸ�rH_� �z���$�r*쟴�Oi�B�!r8�9#��=��[��X��d�mU���2q�˦���1\}�Ed���)P�7%Tw���JU&���@�Q.d�3Hv��{p�e�a��`"��z��I�e�\KQH� Į-H����o7�~Y�C�i�@�����W�����k
Z8(����^�A��S�
=�S	�<_P��W�Zy�,�~/��*�r��JHF��3�be���kѻފ`yH�gUF����sS@�"~G�M-Z�3nF�M�q�^�������]�:t��u,�Tp\cM�.:��d�\E�Pi%�aL�c�ݒ.��Er�56szFwVK���P�>G$ꏮ����a�Ly�n�,��yH��
��X{V����`�*�������:�L�}�cmo�aF�i����@y�o�W�q�I�6�p��/����֜4��൯<L)q�$M��+b�+0&7��~�p�,�7+�&�p�7|୊����`ʠM%� վ�q�T�?���1	� ����G��Yd�q� N]�,�U�,�3�j5b����=4�\��;��:�f� �J�ݏ�f
2[�Y,�:<�� d��c��'{l-z��'�a�|���/&T���0O���ݼ�J,�7��t.��;�0
z?\��RY�Ŵ�:�޸Jy(�ݸwm��fAZSQCƶp�4����MDqj8Z>�(�n�8R�Ҧ�3ǟ�����^xG��.���(�X��"�\���[�f��6J�������´g%�I��j��{w��C�v�2>70�M�a���?�M��.�Lb8��	�f"؈o�6�]V��c�r1N�cP�9R����L�����!�����D��@��*�ԡ�[s	���p��Y�q�|(���C�UĆ�֧�D3u&j�N��V)������	�(�D��*��W��pVJ	;#�\I1������j ��p�{�z��5�`mz�|����(�J)W~���<�)dh��o�A��:�~�V�"��u��s����b�Ӣ�R���Ma�&,k���%U��͢�d����~���X���i�w��Jw�����HBF�=}���NsK��e��Y\2�G���V����|TYDN
�A2�8`ɴ�"ߠs{)���"�:�@]��G��6-�V�S�WE�8�ޘeNidí�ݔ��,;M�j�Y1�=�� �PL�W��xw�	ً]�3B��{r��0X��\�:Z��CL�=�\2�디��\��6+�� �ȡ�8zCH<]���%+,\F�4iP��8V�?z��`!|��K�=$�|��rf�z�#K�fK=��g[]n�8V%	��U�y��)��]I~T����o>��K
t˪�Z֞ s\��\�3�Oh�o���b�
j���:�j������N�����5���=�6qZ���a � @�\y ���P�0Z!`�e��C�6qg��T.uW���=�HpZ���z�QU"��q�I�O��ea��H�i�C��%����E`.v7T�*��r q�X�e�y���{�֎��M_�7Y�Dj�vz���8j���g��\JJ@ɖ�1�'�+mI����_Y̪�n� ��c�B�F�1Q�G������mW�x%XWPd�h��?����s1z��z�t��O�oK�[~���{5'F=���Ƣo�ZM۷l���X�_^Oa����#ԪU>1����.3q��(_�(}�?��$*�T�T��^pj��}�vG_@���o�ۅ�b�q5��SE�K�r��j���7���k9�z��x�#��q82��WLJ���C��6��mp�g�V�a0L�d�J����c\��_j�5��Gw+M8�2d���m'��)"Vx��_ޡ�AQ�Ҩ:�_�aEnT��E�w���A�����cUiS�Ҩ��6��Ex-�� ړ(���J�l0�:���?��^�1:�Q>�^���k�셿<��:IF7��`�uP�+l3��y�%�l���+��l��@���O$��S�V�2}.��P��Y׬�N�'M�~�8�H�J�u^�L:o��bQ�n ��ڀ{���&���Me[���#Zm��3��Il&'S\@x�騂�#�gao����A]�H��fL�I�N���&K.p^�R.K�O�x]�\�g�E�1��`�����>��t��Y4��7nʡd���-��%'�iK��T��d�wχd323ǫ�k7UdtQ�o#F�G[��&'bc��y`t�8&�$��?ɍ|̂՘�a��LFF
��Ӻ�`ϙe��v��B63Wa�k܆��n��������2VOz�jidt�P��(8U���{56Q'�m~�MU�\��
���b(Ly���t�?wM�n�q��u���C#�{����;�yLBϫ�����a�e'ٯ�v��oy�M�i��iq)��@�{Z��o"Mº���b�(� �zҳ**��.�r|�VٴJ|�^l g��	������m|�L>�S�E3��x�;!�)m7�@����!*U��7X�T�PL7%��.��!�>�T{$7�+(����tG_.B5N��c�Ңoݓ)	 ��2Whr����u���it�R3��)"�����@S}�Ԕ��X��N����#T }�<�=�8��㷨��o^K�C��^oz�۞�?�^W�lQ��B��>��˿�̙�2h�}�$$fJ�O�����;�T���e	�4�RՊyl8�|��]��AZ+�����I�V���M8�gO�u�]Q�jHb"�����J��W�m�K�6��*�E=�ot!/[�a�/C�*m�s�H�Zt��e�J`�G�42x���+�#���8�xD�3�;"F�/ %7�!���)��_j�cjξ��.ZY��}�.�Y��/Y7Xr�F�{b+���eÈ��0��|o���y�bn��8%��eNd�g��	9l�;��i�¡9rؑȍnI�oR�����gެ�IL�uĒ��5�����/�.�br���!�����-�E�^u�;p.N ����#L�I��(�7�"AeVu�yF��� O6�]���l��)�5m��i����F|~�R�23-�C9|����il�oUg�̖�᪦z��m��;�"������H�����oS7 ~���u���[����_

zk^��n����]��R�h3��v�Y����j@Yd�t����<"_ӥN{����tJ�����QĩZa�yx�<�>�~� ��I6���2	���M"�=D��ڟ��3��x#z}��PY4!����å�����z�����f����p3�'�`��~������3����ҵ�=ݫ�=��o�w�:=80����A
�N�����UJt��-Qy�Y�,��k�En��j�9��׼��4o^¾����cͤ�,�{W�(���F�c�W�6�*���_�fx��U�ǂ�7��t9�K���f�cرCz��!ݼA8���i�D�����7W�\�K��7x_�+���B�lW���\����P~�-��q��0
v�.�KS(�RR�������98mn�.����ݗ�`� SD���t�S�|�0٤��T��ٞ���Uۯ�����8��M��l^�&[�I���HYwqp9���0R戯�͍�L'j��}�������Q; DiS����nx��EڈH_��OI�-J���D�q2ٛl����*�sX�X��Y��=���6s!#�[~��U*�����B�nT���x���W�I�kh���i��!��4s&�,�ѯV\�/�si6�`�\����sP�8�بH�ӓ�Y>,�Ѽ�Z��a�a[��).��ZJ�p<�����)Y[��I��?��~��}n>��w����70aX4v��)���h���V��H���x�Î]9lwB/�2��1�<�lӦ���V�[���;������4�gV4e;+�X��k�b���+�5���Upѥ�q��F�&ia}�����u#/�����H����^2����͙3�}�ҥ:���p�%ٵ5f��K
���/�B�D�~ې�����p6h�A�sV��.0�t+k��Y�9�d_i�����X3>(I@-"�[��Uy�����ZT.��"�y��4�Ԛ���Q**,9I�r��d�H�|pҥh�m�o[�+e_�q�ԅ������#��U��#�F[ ����{l��/�K\�J]1���6O�P��k�^�����k����<i�mqc�/Ay�M�\p��bޟ���s�!���嬻�����}�Wj�=��%q�\����[f��Rn��~mȿ17�s�:�(�����î�^HIy��Fe�t�Ҥ�p������A�w���R�<�BW���i����AH5'��w%}TBQ,��-��~E�s̤Vc����T�$"�z��@���H�Ɏ |�����ab_�r1M�s
�k^���. �3���� ��������i�]��a�~�5�M8_Qؽ��DK�o3zD�>_��%�1��F�,0�FlP�O7W7X���j�XCEB�{~sJ�dx�[~D�ғ��"�������ha��T��������ފ�S�p��}wjw�ot�v����R�T �9��f�!r9	�~��a���)��r�F|X�=dmz�=���bN��t������}�8dܝ��9|�W�ו�LSTT��[%����`N+��qg����`�;��:����W+�M���i\BT�zlu�赻L��l(!�-��d|�/JB�}�e�Kc�(��<�r<~���#����������}j�䒞Ub��%#�Z4x��!�|��H�3�b�`��}�S(W �D/��fUj�p�:�T�vb������x�6�sn�� 8O��d���Q@':��D���&�gK�����>ࣛ���Ӭ�sٟQ�Rئ}m�]4$��B��� �n:��"�gm�'��w^�,L�f)a�.���^ų�shgBk����q�K�i�!"��I-��BJ^)�RJ��E!λ�ǌ���>����**}r�����@)����]���9@$����{�����dR*c�}���>����`RECKЙ˒��ř���תxDRm1��7�L�u�?u���S%����Ú�PEs�K^fiE�P�RgK�h� L��l z�礢C��Zh�.+�g������Zʍ@�@�0Z/WbN7�X3�V�ڿdt|�oL��=;���ᢺ����2M��=��(��"�\lv]�3���v>�tYNYT��]T�gz6�\�,��1���Ƅ2�1F<����f���d4���\��t��;Z�f�����;�������/u�9��\
о��D����h��\�/���,5�� 0�U%��(▏�������픳I̩> �J�?���;�� ��pW�/Th�3��9��La��w���R��h^�"m��_Ӄ��)ݠ�<�J���Uy�)Uo�	�U�h� ��$e:8�z��0���E 
*�2��&]�m �vʮ�!K��,<����N�s�H�߂���йW��[�N�3�|76Ң��z3NN��_��E�u�"&F)5�b�s)�@9�F�9���b4;5�o4PS�.Zp���ؽ��I�Ui��+Bn�+9gQ�0�w�Ce��Lr���b2���8�9&�~j�ni���;q}����kUʥ��z���E~s�}��C�R �/0�q�'��W�v�_�=JK�m�.���;pg/P�i��!iDh .��$+M��f����!/��&�6=�3i
�MG�Q�[�K�%�t��fvz�#��m�3	]"ف<��io��a-˃4����5���T5���!6��F~o��;���R����},w���j���f�_��pu�h���e��ֿ�sH~څǾ'�����E�0Ц^��r:�byONI�M-��9gN���qV/���+C��[���_�MfC�ܝʲ�eN�����D�{�&�yO��dn����dl�${��OX#������vd�l�����A#�{��0�����u8ҋ�3������2�2����}��������ݽsט�t*r?��0Їy��C�!ۢ��qF��Ɖ�NY�B�ɲ0j�ֆ}�W�ٓi��Ċ�H�5iq,5f�1�<.!�w�� X���Qy7#��|2�Bɨ�{�{�"�� �-�WF��܂<�sN$!��#s¾�n�yo�j'���&���>�3��|S��m�#�W�H5r�b�	������f�-�Ȯt�^��)��f�8[_>-�Hj eL0�>*��B��BCƤ�OjH1���r���c��yʳ��K�Iv�gڅ��q�F��ৢ��zC7����+�T�>����Mb'q�ֿ�Cqǲ���^�2c���.��!�a����ʺ���k��v�300��nh~���0Z���HB% qO�J�T͵��y���C��޴�NZ��c�/�"�Me�RX>LdCc��AR>;'��ͽ�.�ǉ�)�=�t��aĵ���%���6w�K� �z�E�i�׹�+H�>�.h���b6�՗�"0~l�1ڋ�K�Q�!�ۡ+�@�T�H?�S��fwҟ���έ%Av���1��5�-qy��,�5�5M@��o�:&J0L��)f�|�'HQ4Uu1/��0�D�8���L_!�=�>��ؖ��)�k�`?"�?�BO�yܳ�P7�)�^hE2:�z�����=��A�v��"��:K5B��x?ձ�Hb_�#b�-h���/3.+�?����o�aQw)�_15�l��^�Z���EW���H�ڑ�nݍW�}��|b����[ԙ�å 2��lCiv"6U�vC�jr��KI�_F���ie��Ə��\f�R s�3����&H�]��ϴ��h�)y��n�1_H���/�d��k;�l�W�|u��/���xW7￱����W�������ƀ����|���s7R��I�	���X��Z �_[�L#��oZ�ץ��Xs����[?��� W,���uM�A4R��g�j�S_�xw��3�إ����M��J�������apUj�\����yP��]�j,2�j����;���[f�3%���u/I��O�&-�B�;��oJ����Kȩ|XHY�1��L<x �Mv�ZlN����!�~�lk;N��;��ׯf(���[�A=�6�������|X��D����M-��Ͷ�'��Q�i�hzO�C�fA��<]݃��"-�f�}x�^�B�R� L��'�9ڔ��_�zU�Z9��1��RG8�d[6�%�K�0 5Ƒ\�l3@�p�x)��V)����hQ��h�c�Ї3dʄ1�Z8��dĻ�����(���D0'�0�Ps���f�'�q��n~�{8W˪KH牟#?&ol5Sb��\�2�M�����,r��tJ�e��Z'���Qx7b4}"[�,-O)z<�d�F���rI
�9�+m�P׫oZˠ�3�y�~Y(G>�����h�G7����=iPz���D�U��zV�3�٣e@�?�=�����3��<p�8��Ϡ�[o�_��#~�g�I>_����]ͲA?��f�3Q�m=H
X�y�@�B��"�믌m��$���������x$c5fk�b��}��q�p!�����S
�z��������N�����z��TP�}8ٰ;�b�np.,�ş˳���/@�E�]�%e��x}g/�wA�Q|5�`K%@��.fF���
{`,.ac��sƵ���K]��rE夎�����U�_���(��ǔ7) ?ڢCE��	v(߈0$��m�U��P����y+�����H����
���$�=Y��A�w_Y?�g�*���M��!����iN��q3g�o>�/}�qC7�!ĶE9��X$:f<j���@4e����hߞkD"�uM�?J�`ȯ���pK.m�T�&{��{�tz�)�<�|B.)}Va"�����
���F��J|R�p���΃��^��1�����KS[�׻A"��F�]��qL��w�����H�lL �Uw�t�BR�����Gbڵ�
��C�*'Z���e��=|��U!$Ɨ~�ƺ8u���K��:����+�� ���`���z�o���-Å���Њ�]��š�m�Y�T)�:���`T?�����U�\�3�?�A��#t8p����$$ܭ8z,��C�֙��v��� �N�ӥ#�Е��DT�$B��*��
����� ]D8���yXM9ONZSѦ��;�IN����|�z��L..��q	ANɣ�H����+�I/�l�a����;��;�_��_��8���H��G�a��}������Jް�W�{Q��hI��T;Q$� �u��&����: ��;���x�_yGG5��p�\�3�"a�x������R>�_8\�4���ӟ��E����"�Gs�҆��JUT#7x
DN)u�a@�f^Z�:�G����F|�ޝ{��^l�jQ1��R����A����Z��ȁ�yA������CH)���l�q"����>��zS��?���{8k��i�]Z�W�B*y��2���S���J�W{��0����6��� S�2�P^ ������㎹+�x�_����٧(�?�!YG-D�l��9Š]�ζ}@�kp!��/���	1 �\dzy)�t����	{�ǂ��%yE1;�f���>E�ޗ���!_�	<���ɥ�\ب�_̓��H-Tb��Gpd�-��$:p�"8�E�0R��0Z��Y)Д��l�3E!�R��y�yY��=ן��!;��D2�Ҿ~WCkc� 3����U��UV?"�vг1qtI�𨦋�����<iL�6�O��1���s�(ɴGV"��OX�y�2�i����q��^C�b���e��[���I+����u�ȅ�-���X�g�Τ,k��(55ml�U{�2.��s����x�+��Wh�D[h�J�±��l��	e����e�K]�{�i1�up���`Ioy�0��� �qXe}�/3�vҀ3�9���ymF2�̭~�wۍ/�$��$����6�$NRF��$��W:��WSxw//����T/��1��}쓑^�Ƥjh1r�צ�'x���F+��j�����OI�'���T�v��U����E���ŉѣp�.�����醘eT�á�w��d���h��?����w���y��"�r�R�������Z�D�Iu|�ܹ*-�W��$Ҍ}��<�^Tt��\�.�\2�%/b��������EP&ύ�3u���8��S�|1�X�e*�k	b8�Fq�u�@�e�m�7�L���Ts��ī�l?��8�� a5�I�"��Ie鬗>o�|�_(?]C����i�A6�����c�@a8V��L�=�h���@&����t�[b�k���HAlv[dbXV9e|x�:"T������]>�ڰA+��W�l�@-]T�
\'���Mߖ(��r�R	����^Tܒ����� ��[��T(X��N�O��?;T7�����ҷ*&��[�N#����%�䍖Z1�u�.>,sޓVk���Q�x�HA:_K�0����QLV���3����%芳99�[<��[���I��n2��J��9���~(*[��!�#�m~O��]r@�6�gemo�����r�^�=o�ӷ�R�ul���Y�|�h�G1��c���!� ��I�#N,ª ͌��1~�B2���f�rGF��~I�M�`E��~�m�!x3�VH_��.Ǐ�}�|�94�#�dT����'O�c�|2#e신<���W�˒�p�=��t@��\��r�n�Uc)���S�Ɲ-�do�������J�D�#����_8��H�5˻Oe�j�y)��mP%дe�Q,ϔ$���[�!��D:��4����)��[��>���U#����q<�S4]�Ǧ��C�'+,qc��3K�|�%T@d=�@��ȶJ���R��Nn����~k}��ThǕ�(��X2��X�'	��>�R�r�N�o�$�`�(j�P 7��U��oqo?\&RjI��9��=1�z�3(1�j�L�S1���r�f����'�BK�	����{���:ܝ�1Tq��	�T7��'�ߖL�XCCM3�7�����}�5�Lze�Ј��;.H"��%n �.qq����[�RR�l��n�Ќm1���O��p4W��:��}`&���'{������u(z�� �� �܉[�^3f_p����n�щӵD4Z��6��F�D%O��{�E����-��#-e�@O\f�o�ʄ�|�h͒ok�N_Fc��#�s}s.B� iG�&�	��ُRmP���×�.���x>,mܹ��ű�m��1��9�u,�^�=N�������Ѱ����0�ǘ2�Zp�0oP�D����8ѥJ�#by\;#�~&�x���N�G��^���V�l�V�e9�^VX�����X��G�Ɣ���hOǀ�a�<���цub�8�_#�z�@H��{�A�(q�q�ܜH�P�7��V��$I�Qկ�
Y^򼶗W������C�<���'�1Q�_K���	�!�c����� p.jV�D��A�����I�b��2r�M��#@��E�IԿ%,e���BÁk�@�C�k���B�L"�Ǹ�H�!�u�����)��n�"�챍O��d2�%�4�~���Ȭ0���Pس� 
�F3�@@@a����rw�E��Y���k8���U�Mi�B�C�\5+㒅��Bf����@\��.���[.�-��3#�$�Ҽza����U�OK�CG��r*_:a�އx�ү<ȥ
��*�U�Z\`o�Ν��|�Ԩ�ߧ�7ɏ���-�¨�����CAb��'a������0h+5h����iv��f��SU�A����<�RP|Z۹6w��s|�&P�W>t��P���+��Wy楜�bڨ���g���Rg� �r�qdJ��i�:�^]A�ߓ�g�3�@�_��i�#�y�u5cs4�2�0�Gq��BU����<�g4Sr�L���Z����<;9��K�Iv(���w ���1ɡ�b�\���<����x��CPY�ZW5fW[���ꜱ��"@ӱ�t����&:�O���tfF��+̾�*�$ıs��
�<�N���?����4�[�B�Ycl.\Z۔u����mJ�.���a|����Ru,~c��>E��R3KI��2��O{�R���)�j^���e!�w�O��F� ��W�u~����ۜ�vb�]�.�����%�*�o�dܻ�O/<c��!�VDr�U����#t����v���y ?�x��V\Շ?S��5`w�q��LJ�&��9�QiQ�%z�>`A���@4k%�9c������t����4��V���`��x�?S���J@�O�þm�%�L{,=�Ǎal�1�Q��~�������_�H��K Vs=9`Jx�+�PK�yf�>w�m^~i$��M$�h�K�	 �H��`5 ^�7R�ɢ2r�u�Nؿ�E �tN�q56<Q8R	i{Id�7l�>H'ow^�x���J��j]�*%���I���9'�0�\0�W�fڌ~V�˘۵r.�P�Z[��2P��^�5*�L�sv�B?�.�2��˥$�9�]c�/X�dw�[\;�����ZD*1�߃�Mc!٠��9�N��|`��0��%
.q� ���a[��q�o��ȝ���a�mTP�⥗��9�|W�)���{]J���q����[���b��zE���_ŠK�Efw��>�Ƨ� ���"����ȓ�h��<XX��?-SU�?`+��C����a�<X�L��lgk�2�O�S�f�s,�4����͞�>CQ�wYp0���0���}
�#YՊ�DaZ}����&��H�[웏���`���`F���t�mC�H�/$M���^<H�f��=���1` d�Y�����uI|�(���\(�n��갶zT:_sg����҉�4������M]�6&g�ݠ��R:��әsōxDH�P�nN-�A܍D�t�Ӳ�Eui?j��/ʘ7��:vRG��p��[0�T��5��$���O���H,>�#�����շ\^�tiY�ţq,1r��KR)4����S��J��O�]��Q�	�l$�w>��4�`�RR<�_�#p!-h%i9+�p0��=�P�ARW��/�,'���!Iw����JFcS�Y��)�k�t�51ȕ�a<��%�ݣ��tO廩�V�Q�K'=t4GU�= ��������
��$\����Esr�T�|�&�����Ɗ� !(�<����{TKT1J�X:��K��;�9���Tu8[&� ׇ�c��$6")�J�WǮ�9u#��.Š�'=�#z�SE�S"��\�����N^ٜ���o��/j"�cK7tϻ3N]����pc{��y�\�PQ@�x�j�ВX�K��d�bb>��IMP�گ.\V��3�|���O�:ی�|��\�jX���}C&q;�*n�[]�X5c�!̛P�]�g9����~c3��.�#���c�ּg{�j��]����]ʵ_�����On5�H~�-4�"��<z��I�T"�S����8�c�#�#8&^�������_����m�2>�­u������'���� Z`SHK�.7����P�wtBػ��V;���$���T��T�d��܆�&�(�y�x�
��`�3)��M�v���Ϸ
�Z �\$�̖��g�0%��f��[qY�k�R����g����Z�6s8U�u%$c�d�:��b}%D�B��:��{�~��O�d���E��5�S�vu���=���S�,t�d-?p�j�ʫ�o 74� c}֡&�&m���a���/S|Faw"��!��CS�aD��J;��B�Q�#�	@�b�eɄ22�3 GdXJ�9Ĉ�ڈ�|�n�D�˝��?�E��8G�A}AÍ��Cm��T�n�MP��Go�P�U���)�bm�*�c,��q!b��/P�t��i!����FU����{��~�I����U$�<��d��1�XT���O�wf�҈���֗L+�=ca�P+�s 7\�P6���^\���6K��v���K�g��u2p��R?r,|�Dq�Q�J@B���M����,pr��
6-Ðn�y�HCCL����x�!��QD������������jȮ�t�Ȧ�k�B��4��;�e*���jԋ�$��Ѕ�":'����{;��!�<b�/��*� /N״��ۼ=����z"�v�I���],{`���&�,RO�{���������, �I�����e��f���R=.&���o�����	[��Y&JbAo�y*MR�GMb��6�0D����@%�@ÿ,��������e�5;�Nr��%sM�p�~�gik��ߌ�q�j�x#�-�,����`�.1G��PH��M)��+Oc�㗃��%�UR��`��(iY�� $ݏ���:��H�+ه��y�w�eO�����ɀ�c1�@g�^+��C"y�`�p#����]�fH�et�_�h1i"4�x��3�sH������<��H'��A�0zqϛ�
�(�a;] ˖����o�&���mn㓮 �k��:z�������#���Ɔ��(���L|��0�#u�>�$��Mo4"n2fɗ3�B���)�����;���r~h��R /�'�r�<�(��t$_��&�gjC4O���.Iz�B���ܠ�ي��H�x�Q���jC�yy�)�Z�Q�7UK?�����m ��Y�c�O{�(��e�.\�+#<݅�� ̣H�-����t�Oyj�{�R� ��{�E1�S)�խy�Q<� u�E¹��F.�w�ʈ����ܔ�Z�"fJ �?M˱�X�k���V|F^�0Xܸl�KD3q�J�V�}�7N�Ĩp�����B���2Xu�e^:�[.<�n�F��^D����r]nSDn����+�.�#�I�*�`�@�`�5��2�~_�`���U��os+�\Bz��%�@|��RA��]K��W����H�$Ì�珳���ouk"v�8��I�q��∁���� `\L�.p]\9��-�-դ,��w�݀55�3H���ZH1��ge�Ls�U�kإ�=��/�4��eG�_FrR�������˱+<�����>�'�vFF�BW��:s�R�F���W�f��t�v=�8�S�Y�#S��<Q���}?�W�D���W~)
.sG3�/��\�@#W`[��:�@��{0zb�M�n��`�q�zm5 ;�xQ�����_��_;�]�-b��ʵ�I�TA��=j�A)d� ̙�Y��u�2���D)�˳�8B�������A�5�}?Ŝ(�U��C,(��f�h
�2]�aO!�&��ţ��靳'}���� 
��%�oW�w�
�|�H��F8Fj�bۧ���LV?��[/q�����a���h�G���\7R1W|�[⭆���`��Y��}�.I=Wשgs�@������T�������n���Y����d�wc�M���������`�N�P�%g�#�Z�]�!X#z,A@|p\#�,�X?_{�C�|fR�|;�)k7�C(!�k��a��.��d�`�y�A�3���d�
H�!*�G��h�/f��`��M!pͮV��<Ư{UD%�P��^����~))F�H�*���|^�b����{d������˃�y����U�Y����nL��T��v�+�Ü�i�Q�7~�B��ߛ�3���ۺv�G�T�_G��!}��C+�5�����Pg}R�]��h��e"K�?Q<���슠����q�2��Z�C@Q���M1��.5e5A*�@��	_��$�s��+qo�U���5��Yl���z�m�o��a*�7�<�">������9��5�Z|��\nڛ�������lk����+|��cD��B �+B�*!�e������ٕ�P���\�㞗"ֵnÎ#d>�_GS	�r~S�걢�NW�ir�d!A�HӘʛ;�\�h�:�67�S=��	��Q���V���;����D��D׃XM�#q�x5;5dT��N���<�-4 �"(�0mױ�4��,=<1pq;=�9p�����=d���V�����A-�% ����D���J��7�)�a�*�ˌ1�M�2&F5������c�8gAbdd�Ӯ��� 	2μ	$T���g0C�k�53��U[>��N#z��ԙ����f-/���kV�m6H�`C������J� ��g����#m.ɟ�����8a3e��]�F _����U�>9������Fki,;c��-E�՚���"�X�q�3���Q64��,9��Z�4,�p���G­��v�������D���i��޻{���eՎ:�Dt��a�u��
b<��!����I׈(�l��^X�#9�6'&��r����;���!����%�T۶,��1-��$(9���mp�[2����8�o��;�#�Oz4���7$����Zf��@�(�ݔ�ͦW�ꪪ��o�@*Uo��f0]�#�x����F�'1�٪s�<Y>
�0�*�Q��lή��	��\�m����:
��Y~��!�j����/���p
��rK��L��+���}��$W'&���q�Ϩ�ҥ�ƻ� #�荴ā~`�?`C:o���~�L'��	s$�`����'�q�TM�B|�p WBX~B��'�M�^`�`g��V�=��ϡ�0!TmQ��N;H21�I�mg;eaT�Ԧ�}��KLpCN&J��є�T��#)��yn���U$�@ʒ(޷P��ʄ��<��uL�R d�lH;t������V`D���A'G~Ӿ�&�׳�ؤ�,�]�A3]�8�J⅐w��A'8��H�(|y��?5�"���!�fȁ%h �@����d
T��\S8�k'�پ]?�YͶ�ܞ�	(��s�ǰ�\72�`ìǡz.9�ғ�#t��J[��5��$6k��R��{�	�x n*L(]-!�������Z�T�{jz9�A��rc� '�]�"q�O�;n5r�>8���X�
T/�+'����F����ܑ��n���C�6v1�7���g66!����vZ�kAR�H�e�#���3}��C'x�Hwy3h��;����T�Т)�aK�?
�C=�$���v��B	��, �Բt�Rܮ����q�����"gb3�7O�ߊ�0a�<q�z3�;꬀���`�t I����mpD�v��4���F���\Y���sk��;�U�	����b`w���hB�uY��t��糐Lٌ�'Qe7�H�TV��N'x4)5'���Pn������vu���
��n%�f�G���������~�����-t:�<��'W��J�a���xpǓb�VL�4(���'�*!n�h��c~XH�-�.A`��� ��#��U�av�
?���9D��6�n�O�o
�]3H��=MD˾̢�������a�̝M�t��g:�ָ����@�"����F�k݋��2�y+�� ��+{i�N<M*�ݤ�?jW�Rգ��uK_���Jy~��|���h���֟�#���؞��`������c�.#6����*��7��:#�znPO$���E?׃5�����e� ⴚ(lu;��ݕ,y~�%@�U�� W�K�"�W��QD�h[�u!x��TT�=��?p�PF�����*�pR��⬒JM���ĵ+��=���]��pN������eHA-b��ğ�H�{����)J�VJ�;�3�*(�Y���4T����s��@=| �����?���`��(�R��f�1p������<$���	=A�K��/�0��ɋ��BBM;Y�@{��K���6���[S���m��)�mmx��[f#�0}:rO+�V��ɛ|�L��|��SIR�ґ�a0s�J1Zx�R�\0��m�С=�Yf )5d�.�v�qH1[����[���,e��jAM�E�A�`vl�A1�e߇-�]��婺�yD��*s�X�O���u����-�n���B�����w�y��q�Q�Io���%�������n0Q��p������#�VӢ��?7�5�Q󪋟.D%v11��M��^�Jd�Z�3����k���a��)���� �{���=�B\͂����L��k�et:�.�	F�ݏ*p������@��$��.��?��e�E�1���:�´����*SQ0���[��SQ��J"��c�sM�c����#����3��A��Yv���4I�m�|\I�����l��[b��GI�6a���n�Zȯ�
4lUqW�����V�[B_;�^�^�l#o�����.}�>��j>�s\'�{����P��-���%S�̔��hU��Ԩk��sSZ�}�`�d�G~Z��7tk�W��P��n�]����7<e8��O�yZF����`��=������410PQ�>�HOnfLe��:�*�� X��$��
����ȑ��6��V!g{c���cp����^"o�-�$��A�6�$!7�=�����%RC����H�V�;2Of`Y����<V��߀��1������v��ɾ��oz��,��A�����s�&���Aƫ��V�:FqF���kLvŘ%� �*�##2�s���h��U�GE������C�Jʰ&ɼB�W[:u�M0�X��C�ɤ��\�+���v,aLu��ɝ�6A&+G^د�\�)5�+��ʹ�W;������Kթfֿ�)q�|�F(F�;ֳ^ͦ#Z���lAo�Ym��K2�b#��l�W���n��lBTuW�fG�G�����~rŶ�H;�P���ܮ�Â��D ���oK�������[{�G��|��o��jK�r�`5O�W��7�i�JtX���h��K*�����Qind�UۯCg6���j,#7K�:ct l1�r��,�k6"���A�s�ȕev��l�����7_@e��f��׭�${�������b
�_��m��`�f]:|�}�-&�+D�����k����b��_��p怏���/�nB��G�[k�U��,ĩ�I��@k�i�=���l�.�o]��=�?��'��C�Mi�-"^v��V�DR˩(B7v��';��32���!�-yId���\�V��Mq�w&#� 1Ԣn1E��v��RK{��7��瓨p_��Z��cS5�7ƥ��v�zy�j�g+TF�k�	�\;AS�t}&���lq�mޕ��<bH��ۨul���:&��`�&�+uby	_U�h5����w����4��%C�Mw�U�)y0a�S��~�M:�'��^@ץs����R!�_HZ���i�yn��VڟǬL��Gl�-�G9I'G�=ժ J�jـ6����3{�/�p�ۊ�A]ħ���0�+{�3fX����CcmE%�tɧ��n�i�}�k^�ej�7Kuͨ� �O��#�,l���Ēe?otX�_e�|�v\�վ��b��mʹH�X��NϏ (c!-[}h�r���K��NZ�h4���!6�%C��i���a4ج�9T8�}(AM=��Ǌ��(�`�7����XPFܛ�IS����(��l}���p�s�O{���'����
2w��J�R�vL�l�ל�P�4�>d*��Û�?�`�T'e�:��sf4��%�,�xe*��O���%V��m��t��21�f�>�IA��:�	ۛ0�ύԎ�Rṭ�gܪMU�=���Ԩ���n�g�q[(q����q;�h����X��ء�.���X ���a�"�=�A���H?Z���}-_B(6��9�)BUꝈ\I%�i�W5�G�iJ| ��d����4W�_)V_Lo3��;@��8@�ˎ��� �dD��P��u�@�],�=ť(x�aTW�شۙ�l�)��=� �P�A ��=]R���������D7c���Q����VO3��t�% �yJU
��ʪ��f�k(�Bu�W����"�1���͗���n ��jƩ�݄P��ݎx��&��H���cF4;�҈�CB5xF�@zE(CD0,���d�ְz�dhH1"E)XH@Bt)8�n����l,���if{��JZ8�W�\)�qk�@�a}�,��9}�W~�|SR�/4�"	;�N9&Ƞ��4��wd,��l�%Li���`�Y6۬����a� �gN�03��D�}X(kQF�"ߨ���m1�I���T�x�Ԛ}�;+���l��T�w��%=4˖wK (<sh��\�t}�:�.Z��?\N.}7��gCRcJ��0�F���Q 2�bX����xHM�1�ɏ�"ER��~�;5�H_%� 
:g�[g�ȬC`(i�C�pup�P6ps�:pӮ�)O��2 ��v4P΅��{:�#	�3��?�+�?���>�e��D�F��������7�p�;1�{r�ʣ /�2
�J�a<���D�3�:���_2
M�P�y��,�[D�^�Bn����4�� �٘�N/��$��Z�d�U�(�� ��>:��ҥ���(�$,�{��4����ڶ\�K:��H>�-3t[�ohy�=�8����ɕA&�z����6Kg�o7"|	��Ư��q�j
c��V3mo b����q����2pz��u�Znɞ�
|H�w7�g�2�cBks�S�~2���H�n�*�FF�|'�rcCk��8/y�۟��*��x�Ѷ����o~�]�Z��*�6�D�J�$��8�bc��S�n�Ӳ��םh���x���JtڽdӀ�"��<k8����h�Zo~@�K������߃��m�=��?^���������H�ʐ�j��R��&� '�w������T���E�s�TqY�$t]�J��o*��*
�74��^M Q��z
u6�S1՟�A�A��cS����<�"���Hn	�^����pS���c�ms��qʿ���VԾXҦJ	�M_ /ej �m�7���Uս��cY���9�8u*h��W�M�,�����	7v����P�2L'J5>V���������������=P/a~���ɤ�����9��w�wz^��h���s��VO��(c5x�:��
RYl�
Ͽ�q��z���@��f~�n5�$�هs����<� ��.}vݙǮ��R�:A�?�Ğj��0vH�����Y�*���v:�8^2��qt�����L��K��P�u���YxV��+7c�p��wc��:�t�]y�m�acf�-Ok�
MË��E����Gnf;�x�©+\l�O�^f݇��5(ku�B*��c��~YT��R����-UVo��)��:r�L������p�v2��^Z}&�=T�1���q�|j�_b|6&k̀$���Y�{���0�ލlm�ɹ��.�ҷo��
T<��y����HR:p��a���R�a��	p��׌��[j��^�����%�M�ծ������NB��ؕ,8���Ԛ � e� <-�O�w��BY֡*�����6������g�I�����	��J���j���Ҧ)�;t�5Z����Quލ�9}}#�`�m�D��9`ª��d��f�]?�pI�l ������ڞ����cѫB��wT��$��z�A��L�x`(-Gv��q���k�gԤ#��5>
!\�ו�Kbm>�"~:ZDAW&5����R1��a���&Op��W}��|��Av��Q�H�2�����Xź1p<�(m���΃vR�B�z�׌�YI����	��a�I�6���g�t�I�O�k�?n9�*^pQ��p��G\�n?>&�奇��L�|�	SI��������bSӦ�y�:
��0��,�X�zW�X�0�3b���I<Ys�%D�ɀ�����S8���Li���!Y���O�_�y������F�J�[S%F�����R �M�<A�N�c���~ڵY��e�/!���M�3�sV��}���O�s&eZ7�F�sWv$:�r�����6�0$ؽ��Xlg]��m��ڿq����z���q�e��*r��\쭺
��ռ�^e�-/(�a$��۬�r��9�6�+="�%��e*�s̳N��8ws ��tLa⽨����o��5�@�e��锝�g8�wʦ�v\�����u?"x������pJ\YM�6Y�M/X�$`��5֤��7]�OW�h��G���Նi���"+�]� �Da���|R	}��sp��o�QmYu���M�aV� r���?ڸz����=��&��b�&�.s�2�&��7��1B��!�v�GY鐸-��h�7xdVx�c[xf���@�>�˄�NL��Mb!&�6�(���U�d����t��ؘ9``\�a7x�Oy��'�+-�&�m�$���v�i��Q�t��[u�U�s0"��9G���D���ߙ8)c�;��Ô��lJb���� �s��~�!��!���gt�P.�&��g�^#��x��qKd�PW�*��'��������6e�ߵ�d�$�u}V���D@�zf4������ �&�prs��d��0��y3�
{=�?%_? M6�j֫^"��b�����6�)�D;}���1���M8�+��}�����T���J�e��|�By�I�Վ9�1�p�	�Wr^i|eU�u�()Ve�zv@!#�h�݂�]pd�3#$�欴��=��/j���0JԨ5-,�;��a3��E���O���@�[�x ��}$���3����h�_�"��hxܴ/_�8�\�b�/.N�#�D%�zlp��<�{1Uf��G�[ޠi
`�����&j����6GHK�|'�`E����v��~�%gK�8���%����4�V��S��ˬ�a I�I�AmhRU�@�MQ�/�B4&��5i���1�lYե�(ox@�[��~E�%���}����m����� y��g�FF�8P�����S\�d����`�h���ѐ��?t���p ``N݅w�2�
j갛w�1��5_�Im[�Ba��wv��©�.��{�WBk��
��uHx��XI+�~�]݀�6��#HfNd����::�� ��[f�@�U�IA(����9s��6u���o	^Z�p9�m��;�%"�
vw�,� q�?� �m�p�:8��[󇐓��7r0��MW,������#�Qy/�iǝ�D�V`|y�>i<:�ng��sm���Vc�$� W��c
�T5_���Q6�"tK�ݿ��+�K�����,?q\ʎ�$D;=��:���ׯS_pH���@�Ycx-����%�4�3]FdI��쏄�yܸȢu��8�+�>��:?N�֧�0�X���W����;'3#_���FC�̾@��%$����Y?}BH�d���"�����¬밼О�KP�,;�f���"I|z�g��,���ŠPV�k/.��Z�1ȾX]z=l��s��G�M-�������K3g�B��鍯_�@D27��Vv�v�B&��I����+�&SY�\���ec<*���
�)����;�n�!������t0�u��q�N@"������~]w�����q	��'�[���>ʧ'�$٦�u��jʈu�ꕢ�pZ�K������v�w��+���X4M���+Or��l�t:�W}�f�zj��Hh�{̾A0ze������K�cE��D6�t	���U���@N�c!���d1���CN�Y[����ecD���mz��<��Sp���<l@,Ա]Chg{� /�u\�U:S�.(�K��6��<�C�� �r5��i$I�Y�$�p��VE^�v\e�{�DQ*3�7�s�������-n�I~������^�J{��.�q�>d��/ޢ� ��3YJ�$%���!�%��^�ʘU�	-�<F�⒧*���䈙�<U#���<��aE�������?ѯ:�]M���xk��i=�O�_�ۙ~�@���ks"F��F=�.�l�V!������U!޿"g|
/��(�:��1*��:�ln�q.^X�6"Eb��O��,�P���w�p�v��?9�2�D���(}m�ҟ5<����v�3ˎ�wһ���)"7 !�͜mZT3[��,'�؁�3��ё�X���2���/��/H���KX��,��p�8yBh7|�����4o���6����M��
���AH�c&F(�����,f&�3=/�L@�ȝ��X��,$��D��eHsvEo�/:�k��΃���q�f�6�Vj~k���?]iu}��lf��]s)T���'�m5Z�*�0���;��
����4��x6�8���J ��Hi��#�r�]����/��������~Y��I�>��N��ﰟ���چ�%M,���K��=�(с��� ��XҼ��'Z(��WCM,_��B��lpg$ӈ�: Q{i?�<��Vwє�(̟jq
�d����( �@ }��(���r�M�X�U���=��ę�e�s���H�n���� �9���V�K���l�^&�si��}�hU��spX�o�	J8���
�ٶ�؎D�}9�3�$�^�L��lKV]�/<�-�g_{o��]W^tg�c�g*N�4���a��qϒ9T�)���jO��=�D�b��-i�w! �J��g��mG�.��`I_�c;����dzH�Z�{9�oF�&T�!0��W|(8R�@=ERG�TT�:5�22IJ�Haz��W�U㤶�})�vE�OU��p�3h�G9��
2y�-���a%�K�5�]8H�(��"��FgR�^�厂jD�F���JW��v�l\"VX���V=K`����e�H�b0>����P�yS;)��u����?2`$su��H���i�������54��)9��+�;M�>�?G��T2E�I�uS��yZsFa@��XLY���v�]�:��}�p�r�;���n�|���%�E�N
�v	��ŰG��2R�ZD`��
�"��3�Q�� ǖ��{�
H!OS�	����Ʊ���`>#����v�M�`P��L��$Y����B��-����}��#���6��BS��a�L�TY7\U`��9a�#���wQ���BMfX�V�$`�&	��B���k���ZO�2���8�?:�Uj>��Eg���]�p�_.�Ԫ�KtL�P��rrR9�k.�uF��R�e~�T���jK�z��� �hSl�7��c�����y�'*� z�j���@�qs@�ဉ��t~���[s����z�����0����u(Kd�k�U(�m��0:N7YU�Yx2~����b3|3F���T��,�hė�`�"YzM:Ӎ�=m'pssC�J�+*;���Ma:d�8�)��G9�`~��6��V�[�k���T,]�e#�
��\iY��A�*�)4�,ݰ|II��|�a���4�q�T��ZMO6p}\�\���������X��6w�����L_�z7��t8�6D���/餢�iG��ڪ��|�����n�P;�[��H�R`F������mp����HyyzqÂ锘;�g-?�qRh�x�GN�>3f���\���=G���gI+*HA�#��+8h&�{�3�j�492����J#@���]HK�N��s�kH"��G���(��1<�y5wc�n�����DL�R�4����j�ƫ�NL�F�?������^L��"J�0D�B��k����h�D��*]�M��߅��䆍d�Ӟ����t.Ykk�V���h�|�u��%UC��>=���L~{��p�XF�m;)������z�����iZ�mcx6�1{��d��"�m� �npv�[�d7ٲz�!�G:k��@C���ՙ����������)�zYw�x�9k+A�a�m���΂Ѩ@��ͨ�9c
����Ak�ٵ�-���pCq^�[x�%�[����Gai,:)�t�bm]��x�O(#W���0�!M)״?v�y��p$�M˟�]�;4�}�Q��V��@v	�,|�ޓb$�I���/5HK8��1\�_)������:�f�yo��&�1m<2���<�9(x>~߂7���;��lw&�]f�j�ٙp�d��Kz�3�l�ٻ��S��𲵯O���9W�}4�����󎟂!�b/���*�_��
l����fѱ��A�`�cF�ۙ�J��)�U*C&� ��tj����H���2�hP������R����Y�d��"#�FVo��$��|������i�Fv�'�edp.� D�察E��a����A�Jj�Y�w��d:�����2u���欥{���iڈT5a4����RoCGl"M��Z��|!�J���Sn9�C�5����n�K,�r��c#q�b]7=�Ȯ���_��l�=˿�Ң�P3U���]�by5I��>؄���;Qt*7�*Q)-�DSg���ӍC�`1�̐+Ȕvz��LK�j�uV*�6��͟�ٚI���V�j�u#�b	z�����j��≎��}st�9��+��8@>LZ�,�]=�~��:�ȍPQ�xnc��;e�$\�H�g�K^N�E�ez�bԄ	�Ԋh��*$c%~��v�%(��m{ޱ�k��<KvǞ�h�d�K������w����4I�K������	�cqf�v�	DW���S�r#Z}MQ�7E#- *@OS!o!�Q�>`�8"���1#�����*FiM��`.n��*�4G{�G�wm��k��������<c^�נ��w���|�7���V`9㪞'H��\+�`�E巽��nB+��5N���C9]fuͧ���0v��\�f��k����^���ױ�<N�icxM�|} ������|r��)�)i���
��*��*�Ok����Q�q�-���$z��/�<9��y셌�3�X��#)Y���U���t��P��� WLH�ZV�Ūi�8KI�-2���<c_E1����_��w'�-A\K� Uk%�� Mmٞ]$�0ʀE(UN�
e��qa6&D��J���sBPK�dr�h�?^LW-�wzn�6���G�C�CU��>��Q��8�vb��k�MX�q�en�%T)S�������x�I�[*֛!���j'�d�_B��,��k�'x����ud�~��K�Z�W0���|V[b�wp�RV0{��$7'�6ְcf	���]Z�E�9��E�r_{7x��Ǟu!�j�_0��ּ)J����_����"�G>^ӺT����H�,U�6�i�VytQ�|q@��_2q@f�:3ҵo(�7P�z�)s�Ī&3�
� X/�����ׅ�Q��G�%1��BX�D�~J%�i	/«����i���LL��+��r����g���FU�=�ac�4���0����FUȘ��,H^ߍ.3"�����RJ��E��9� |uk���/j�����Y�o��?M\��m��9�xc�Nw��N���S�`��/Ğm&�ĭ��Z=�)t�b�G�fr�9H�*-� ��9GV��{�E)�"jh@t���2�'s��)`�Z�F���?�T���*����,�~zB��3�n~r ��N)�A&���\���$�ib��nsfב8i!W��f$p ?�;���ѕ���V�,���R��uy~�\��Ji8F�H�#�"6���:����GV�ͻ��-J�/�`*yO�8�x3m#Kj&B�R�{"{A���)$v�(�si��
��JЧ��_�Ex��"�߇K!t�~+V>��pD.����3��'SA^IVE %�M/M�7��b0��ݯ{J�F�?����`q��_�?:��\�UC�,h�u�����b�F�!�أY�`��V�,l� ���h��*6���e� b�JB�B� 1C����]����\�. �
ob�Ԓ�N���mq�Vv�/ޥSXˏ���2�(m�kƛ�0$�U�󞘈�c�O����\:>��,l���E3~c� 5�H%��q"���K����.� pd�`_�}�d���4��k�K��7 ��"��ߏ+s?��֢�L
�C6��K�՝%�ɍ&e��
+9�-�V'��9u�l�<x�d��e��cx�	�U~?��9��i�>4�Ϊ)�C���oAV���?Ɉ7S^F/�Ǟu�����+��Ph��˝e����}!�ֱT�� R�q�+�sIt����Uߟ��y�"��^č�=Ep�����MfDt�j��hW�	�Ny�8�7��ؠW^R1�(U�m�C�mQ脻-�������+������=%1�ѿE��P+(����%�^fTVX���^�1"�U/	V�,�q�s��%O��`24��%,�(��/�N��nxg�vTņ���n�z���x�㻪��0t-�mz�*)X�8=Թ�=��ZGҜ���{�ɴ�UI�r����h�R�Q���Va���@��Ҕ�[��1�Y��1z�	��ſ����8cdX;�hdxΌH�l����OԺ7��C�ٛf|�Q)߶3�E�*귆y'�v�_)���c���]Ӏ�(��#@j�v��,����r׼�>�Yn�9�)��?�5��0N��Qf�s-S�Ϳ%���M�D5�N���W3Q��v�y1�m�o�II!�v$0�҃�ia�h<A3��ҿ�wԮ_��{mXp5,#�Y��ޔ�!mz
Y3�c�Y:�`TyT2��~��̺P`Է�Vcۧ��Sq������fݒ�,��'uW��L���>6&[A��yHKS�X*�h��^�iso?P`7�[�A��X����7Xy��&+{&e�B���1�#|�2��m�O�S�/�@�̏
��5���� �����oA���QL[7ʼ��ӈ�Kb�3Ɯ��)|��`�œ�Ȓ��DUܾa��^�����Cp`�d+X!�܌����T��
�h���ٱT�H*τs���ܿ�?�-]7G������l�@�,JT�?�v��L��J�������ɥ$��۽S��S�̶� �ر}���V@#�2��E�B����'�)�
J�ŗC�00�I�t��i�a5��L� �����eUT:���A�d�R"���3���O�
&E�x�$��S�K��\,�Q<h@U8���?�N��(�X�/:�~�4��Y�Ǝ�s�׃n!��u��}���sr�K�Ep���7��ҋ���1E5��j�?1 �Phl��n���r�C6���'e��Sej(�y�-p4��#��S�Q=/����8״U�fc����##+�,�I1�q�Fsx���hb���K
_
~��뗹����a�d�샬 ��|��;�1�}v'0-|r���&`�;b����!Q�d��2������(G=�=���DĔ:r�s��y�-7m.!6v�_z^����;�4?֓f�P���"�8uF����6��8���Ret�n7<d.�XT�����DEK��=����-R2��G�E��R�F���pA�R���kWl>�m�� D.?jUY`���������!dN�n��m'�~�2+��v���<�y�Z����+#Z�4?���j;�����#RC��������4b1�J� ��;�ض�E�@���S ��R�� ��	x���������ӋEaTR��I�^[���|Z�4$?��k����;�;@`C���M������`w�3nW���M;Iژ�h\Jw�̈M7ՖeU�J�0f�!*�U���`۰��dl�rWG���^�K/���+�t����u�8��(��튚D�@�������|kgdU��;f����TJ�[�Z�~�"q�0/9� �=k���X�-�K�)�� ��4�m؍�H��z���r)��*R㎮������ �h �/�k<�3�Ab�����ckk�%[��@hD��,��a�[u3�<o�yWb��7��B�؟��H��\p�m#2���X�,�����%ӕP9c=]w.»O��޷���Z�M �)?��N�X�1����8J��_��b;F�dQ�1�MO�C�d�\�Ij�S?�䵹rF�%�S��[�<^�t�&��[˪��"ai�;�׍��,6Y�ZiH���z��%ӧ��Z�]UOp�����U�X8oB��:��������ζޙ���E���[�� &�J�A�H)�� 9�rm2���Et?�� �9S{�GԐ�i���	2��	]�f(������7�.�@�&�L���oXC�j���
%< Ԣp�΍ulg3����:F�#b�4�����\�P����E�n~���|yu�eC,�fф)�T�f�H=W���Ya�M¹	�� �1	C@�%�udv��H-�L�8K�y�����2��]��.����4�!�Wƈ;�AD-����T�ݕPf{���=�_x��G�Upg�� ZNa�����t�4�o��=� �Ko�K����W��։#᎘y�+�8�0�P���qn������������#�7܈wq��y��B�r���� k��$B��#�G%#�I*��!�Uh���b)e���t#<�j鰁:�;��|:F�BC�9���O`���^F�g�����j-�ݰhZ��َ�����.��ڼ���$���F�D|�ps���<݉��{S�E=��D�͆/s�Xlm\��1pxU_�޷��63-���Fm1�Ų�B�DVCShCF��+0�����Zein��ؖeuDcg9`xéf���.�#�+KF�}6l��|��,���˫��-P�_�Ȣ���N�1������L��C�
�eψ7氘�8Wi���:7�PHw%�{~5��H	b��8rðGsSS�p�5�>%�υ0x[���GH�A���
|��\<���Ѥ
O�2�[����Kd���N��F~KJ��o&�h���5��G+��	T�(靛��׆`� ���o3��H�_8w쒆{�� �(|uqd�9�?�!�O�R!ܱ>Z�s�RI�\��%4nmK=�]�����ad�.�a0�V�L)s�Nh�e+�����!>t�`�e斎�!���9Y����*4�~�(��ע��*F��w6��R?�P��VZ�fF�_Ť�	���O��3���;��lw�A��i�@���è�.-�lDÑ�\�R:�ׇ��n�!>ܗ��._y྾D�ҵ���=�y���ť�+���
dk�fm�j��"�|��,�I���z-�Q�T+���H\�5emj����ꃶ7��ƞ�0��@� 2N�0-�{H�p�m�y��f62z`S�~�H]K
w��α����r�a��y�Z��Ra���b���h�~d�՝N�Π�2�{�id���f[�0�yc���%=إk9M�y�A��BF�8�"��P���2�N@�#n*�i]&���m��jRJ/��Aqan�L�5�f�F� G�z��h��Tm���Az([�\�e�yYߡ��<�6u��|����Kӭ�hNU.��F4}v���/ۦR��ϝ�8j�G�Db0Y��Roh6���@;�s�gאeǌt�}~�4���=�])8�g�w8���0 o��ߪyO���
�i��L�y�7De���p)�ǃ���a[���#Qy��'cǂC���Vj"	؈$G窮X禣�g��Ȧ�aMd�M�|�$I���CZ��w-�� bQ,1����NwVCcg�K��� Q��ui�r���uwǧ�i�����T�����+wo�-�3��8�2@X8%�j<G��'W����>&uiF����X�LYP�G;0iS������hAT�>%�_�?����HC��:I��pCB�љR�PǬ����)�1��7u�<�������-'{�@]��2��hWΡK$C���Տmf(�������ҝc��A-d� �󵄿�6|�������ֽ6�@SRȧ��8�)F��qL��S��[�`�y1�Qg����`��ˈ6鴍{e���p����B�{pKf�����M���=&�~t��Ƿ������=l��D^C�n�I�f��G����Y�#o�|�oĕN��`�k�`�g��{�?@��`�t�0��6������?|د��7E�;��.���I��f�>�@�ny���-��.�L #��i�Q���z=F�P�[B��/�[��t��� �4{H���<�]�Bx��>
Ř��$u>�O(�£���pMUs��Bv�N	���OV�돾�(� �l"����=�x��Y����#��1O�Vi���T����L���S0[�GMCJkW���w�N; ��̎8Y0���[��
��y.C�k劗^8��5�q/A�toZ�o7��^qڻ������r�w�wZsȥ���Eѻ������~�� N��XK|2�&;�:��	)�ɸ$�����L��I�?,0�L�?>�-����������m_ΊO�pc��*$đ�qW?������&	���I�-�^O(I���Ǟ�x� ���$�=)�2��B��W)J"_�*�f L;	��l�n�\ԍ}H0�*�xr׷E�Zn�<Ġ�mi�Z$,�ƆҼ�>_�䰕ќ�	m�I�U*F��M[t�u�S��	�YD"�\%�d��Bb�	�����ۤdAE��������'O�Ll��M���p'}ϣ��3� ���'��>╌>M�=`z_��LH�f?[�H��a�"������(��ͫvg]�B�}mo��#5~�@�/M���V�g��dm���_�%_�'���>E�r)A�}��"����m�o��A��ud���6Y��Q���mMi�8��c\!�o����'Y�j��n��s�5��{y��#��)+<�&'kT�v/� �$vw~�-&��R��3�<�]���8���*G@���;�����7��o�<�`'f����8,Ou�,�"����b Lh�J�,b�J�R�����T�B�zS��]��$�D��ϒp���,|��(�e�Ғ���F����*�+Ow�w��9mWJ��G�1q>E�^��XF1�ONWz����68E9���3�LmVnw�Z?��$�i^(ٜ9W�<�řZ���M��Y�]�6"�[�F���4�k���}�>f��9��t�'�u�r���7��H���U���u\��.aG}xh��)5�Sz41����J���ds���r��2X��!��QH�}���M��K��z�Z��T8���m>o��)X�<Q�đ >whV���/�,��@�dתX��´!��N���.�E�x�F(A�h��g�������1�	�ǌ��YHr�`$��E�1_b1
-倀9Ͱ��n8��j���-�W��;I!��o����CeZf��r�	Cv b��_� Ср�:g�~��������_p�-�&�0���ɾ��6�/U�o��=�� x�Bz��ۻ�\�v_e����I�(>e�����C{T��!��$}T�6�3]��B�9���䯤n���G)�	��A8��|���
*P��v=PD�M�9e�!L�}���b=Zw�����-^����.����ǌS��	o�ӇL�XYT�g����]~&I��ڬ��Rlׂv��L��(a-�4�a	�H*�������Ix���I����7d_2!����#hU9]�M	�C��$c�o��y�S0�8��ʍ�{�q�҈
��ʇ�N�d��vU���4�C����ukiT�xɱp�iDKc���2Tc�J��r���uhsWʚ��9Ǽ��k���k"o����;�*�c6���-����H��������/e"87���}qʫ���)d,v5�fWtUE(ƀy.k�����^Q0�ԏ��͢G���!��&�.�� ��	�)�C� iz.�k�d/�+T�<KY�<Q���cvVsj��W�vt�/����4���L�ן���3�u�~����a�F�\N��򺊖�š����ؾhe�?-�z��3��M'��9��pq���AbF���`�l;�����ʧ��"I���O*�^��:6e+�/�ߣ�ܳ �|�t%��b�h��Cӧx��n�WY쾂��X����gH��ۄ>�s��?�6yBz��#�L�d-'e��2���sK0�p\X�ۖU`����
�`��煽��Z�v��c5�q%bM|�va�d��qR=U_�&�uI9X<{�k�Q��'��1?)�H�����s�"�2�\$�VU��a��zk|��X� n@д! ȱ����M�;�Į�ʼXŔU�3i1�[�4e��t����s����E���|������zR˺
pG�߮\���[Z(���&�y�r�PG�\Ħ0�O����;�@�=@s�.^Y��:^H�q���=�?Rǣ�wĥ�rU�D
�_�Ϸ��	����+�ve�[�>Γr�84���|�B� ��K�����G���9�������_A��`�MzMYʻz�Uғ�;"sV��(:�u;7�ys��q���s�J2�EV������k����n'��|�t<Q'���V胳�G��:%4=�ef!jMYa���@�k�{ �O��0��f����� j}�#C�s��3(�۱ J�zM���H���\R��>��P>*��{�ؚ�{k6l��i��2I��)5'郱��(��?���uXZ߇9>Ǜ- +��Toou�'N�� &���(p�/f��&d�jfEbMY-s���ċal2i��i��S�겊���n�.��ܯ6�t�Pʪ*SA��Z��o��,�]�J56!O��p��W�i����:�Z�(��pO<>����&cxnp�����]����v�l5�qh0���l���FN��&K����PȝA6���\���"�D)yu�.�$�~�_���֘[�C�0f��X�IA9�C/��tQ�5jcR.'ǚ�`�#��9U�%��DO[ ���-X8���Ew\9V	�DԔ�5iK��� ����,��xm�5�u���j0(��U��\a���^�Y��H5�@���:�T$^�ܢށsFTW�1	����Αq�(2�fО^q�>t�.��daw�.����Qh0����d�~=��u�ϫ
a6�SD')�¤��c�4��W��Uk�x5�y��Ӫ�>j�����<�O�� /�kX���َѦ=ꙥ��3[�~�A��#I9������^��;*��I �p��䃎�����ġA!1����5'	���VP�#���ϚFtlq�� �u����y�6% �gI;g�A�Od��7o�_�!A(1�b2S"����
�xnzm�`	�(5����h�4�a��Z%��W\���}o�, ;o�LNO��/0�]��tq��@���6n;ga�Z5Y4-�:�	�!mI�A<��������cC�t�G�.�'w��^���ٹP��3f��'�d���7����4��c�ѱ���Go%׵\g�"VN�0��)��*�lG���F�<m3�Q��X�
Z�<q*����G/�1E��p=�ZA��0���8Q!� ��25���R�f ���9�ڟ����g}���U$̃�Xih��A�{h�M�������y0wB�&}L�?U��UtUZ�e�ۛf������v������ ���(�Hb���_9��{������̂��y+B���p��a�2*�Fv�tN���8���{^H9�(�7��3z�z�DP�`h�������K
A������v:��P�:�b��j���bB1$�P��f�4]��AZU��a��<�-�f��E=��I��mec2����	�b$8<�fu�.�(�%��� ��ȹ�Ս\�#��v>�2���b��D��Jnx�d�O�1��u|^E�%.S]�[�v�b���Ul��S5�E\�SHd>��P/%M�c5���B�Y0�,(	�?���~E��Q��܁����Mp�����]��:Ӊ4�Λ
0�忆���	ج����k4���{/m���qٸ�OW���Um��fJ�xZ��Ŕ�2ԃ��c#��Tm|X�·]����|�]Q�z��r"k��xױ�iy]�t�T�u�!r���|�[�B5I��=A �~���9i#�p%�ju��5$��+d�sf���o%�1]r��I^�9h��<l�t	��?c�`�3r�=<�]�p���<�7�!��߹Z�R�H ^���A�1YLv��t����*� n8ۏ�G)��t���q�2E
g�����U�UE%;��Ŗ��^����o��Yf���$�cx�w��il�`�gb����)s��㚬@bbfļk
�¨���o Wg�Lݱ4ٯé�׉.�6�|�d��Ү��H/�A���� ��z֐�o����٨+0���y �)|��M��%/��5����%��^��N��+�`�k�r��]����??��aU%VbH��N�wN|�Ϋ�����f'�Y���p�L��Z�_�Z4��]���S�_���!�[P�83��E��o�yI��U(�h��z�Jc����q�TF��%�b[F����i�HL�g����-�`sm�ԉ�9��<C�ݾ��O���� �;���+uǎ{�*�@�3Z	#%r��.�|f3��O{��!t���}����d���/>e�C�E���ߺ+�'�>�
c�����9<%���O�]���q�;l�9!��D��~ta5Ұ�b��)�X�ݡ����
�G�.��k��Y"͎��'k�ѩIՉ�=r��[?�5]]F�����h4J |\�c{����X2����og4�ǃ.?���vq[�7^ʻ�[� ��ѵ���kwglb�mnr�gW_���l��̤���4�jn��^�X��*{��epn��Q���9E��7��2x~zj�h�ͣ�4���,x��շQ-r�]C�#��(�U��:��51h�M)l"� ���mm���$So�^��:P��~�l���m�0�%��F��g6����{_�D̀%~$�ة2�R7EH"�Cy[��W���<�����ܱ�6״#��$���CYT�;�L�,��6vJλ�Sg�X8�TM��1��}�I�!>N|l�L+��r��+�TS�w��J� ��U�:��O 3��|^w��S���\��ۯ�@�-�Pu`Y��r�X��t�xy��QBGC���	iA�7�n�� s��^pds1l�r��܎���4z1�L��a����ת35�55� ��VWtN�7gϞ[{~#1D���c�:W�BCZ*y�����c��h��Zp�P7�	2rގ��m:'O�l���+t���r����A���t�08�^\���YI�
�6��ET=Ȗ����0�ygF�	d/��ue�⨄������0Q���[��n<`q�mʥļ���vG�Dz��2r��ʼ],��?$� �Qj�ID�u7~�ۚ��n�M�	���e&��`���n�2~�y�@��2���O�f��N�l[�"�h�J\ ��q��ޕѷ��"���Cs9�z:���9C��(���Lt�?w����Q��gs�	pa��:���-أ>��������V�?�3Ӷ����i:*v����:h�q�t�g�cΤ��Hcd�d��V��~F/�DeJ�MUF�V4�wK���`i�:��y�~���\�R�;����@�¢�~6X�3yS�Xc>+ʇ�/0Mu�z@E�����c��?�졵˙be��ẓ�� Kދ��g
a$_��o�1|�5+T�
_�u]EZ���Y�^�{�?A�G���ȝt���N C�O�>�����2�=�����!�Q�l��|;m�r,%��/ʔy�B;�X�5�Z��M�:�4��6k2��T2?�v됍��%���C[3��,s����@0�p�oi��=�P߉��G�u	\3�5�hP�j��f}IX$&/�ힱ�.�(}`I��<���4�93n���D�l��Wu�u����oZ�oW�Ac�6#�n���Ϟy��t
�D1w�[%O5�Gkx�J��V�U�ܕ��UQ������ T0����+qO�?p��Ny�u�5 J�E�9�����"=����ڈT��됖��8���+&t��-O ��f�kr$�� ۃj�#22i|"�ς�n��IUͧ�̾�ۓ�����9�T�9���|etq=�+�D^!]b�VZ��2w�b�i?���:*DzߌȠs�(��Az9���}�1�^!U;l�j�f�Q }��)�^ eǻ��1y5n�v�y2�13�@&��SEjV��M��;�"��|���)�y�lIW��aГ�s��fv�0 ���ߗ�9��GZԠ��B�m�����S58]�1�D)���J�_1��`G��b�Ԧ�]�����f䍟6��g<�i?+�>`��He��hܚ|�� !$�to�ʛ��,�9�w� pM�z�J�:����x%��3+�����/sCj__o1����j�z��J��,�ݖYa/ֵ1�>���zdcN�*Jݵ��X��o���"e���<�N�й�.?��X���I�r��+@@٬�x�F��X�����#���mMTKn��e��$��f�PaE�ep�Y2�K��$�Ws�f� ��ҋ��}�����>�QX��=K�m��'�F<���+��~k�ĭ]5*���o�Gp�Ι��i�vޠpf�����]�V�&�ք˾\�����K��ٷ��`D��v�kY���fS�0�7Ǵ�<p��7�b\����l�"|~�I�j��!MJ)Ӈ���';�ߠ6[����8�t����!*B��+ԲY�K�����񋅭�;١��=Q�w1f!��x�5� ~�����lőU��\J��+�\�5�N���@� W���S�V���Y�S�2�ͩQ���"����/�E R~��=n�EJrKN���:	�Ѯ|^@�	�$iӏ����6l���Q+��9n���;m��3 �g&k�P��(��h�<G�|�V��:���	���6�,{���?��T�3�7ĸ/F�L��
3�%����4CM�zx���=�����������u#�TH�D脇Qt�O`Vg�%�:7�F�k�i��s���q�a� ��5�PE�R2���#F�TVU��WYO�*�j��� B3��L�J�{�>���qH,Rş�~ b�b���ؓ|Y+��IEF�2v�������T��}�iݙ�7h�=8�
E�c
A88��6eX�]4�>( �8e�����C�K��f¥`�)1��!���޾�S��lP�]�P��c)�e��0���`(�-�`7�[w�uwx{�n=���̙��TXS�i�����<�3����&��L����[�O� \e�n&p�q4:/���P8@!<��8����>4C�%�%�����k��4&ce�<�kN-q��s��$�,A6��Ґ4 )ŗ/{��4�	*�}��O��
���f�/�܏��5�,�b����g�SX���<��ur�����(m95R�7t�p���.
V��K�^��<�˱�Gny?��#^�.=Cz2�Zi;��h���&��(S�Ɠ�e4���F�e����1��b�NjW��V�5�p5F7�	b� Ȟ��7 >����ǽ݆��OH̛f>�\;����<�?��N0�y�5}��5f��,ѹ��"~�H,���-e�I��U��K�T��.&�hOk���XϤ�`b�D%����z<����[����E�s�n�SŽ���&O(���O�3�h��~]!oJ�>�#�co��f�՛"5�;iQ!4M�a,Ő�*Aޞ�'@�Rқ�*r�~�av�Y�c�x^��x
[�v��,�m�xfػ_"S������<��_��Eޏ�y0I�<�>��5��D�cDX�+0߂�۫�	���9�z8֋��U��O�{Xc�d���$B���)u�N�k���+��PVڭ�Ӛ����Vn>r�-�5m�ڤ�]3��PƼ`��v^�`D� ����]�&,���s��Id�G�!R�%���������)@�n����oxQ����n�Z�'��i�J&Z�6S� ���Ux�S:i�<����	x�@S���&��y��L���-!�W��S(!�[!�Al�6o�"?�xZ�,g���U�wtt�O�ECad�����*!eɃK�R���	�c�d>9o�AV�(��/ѓ���.������9Zw�h0{������T6�A[�^S����m5��/l�즂4qf4k�g.��{@�^�cѻ���$w�O+Z1^޵����.�YH����H��r&cS"� o:�-`�Y�A�9W������7P�����I-�<�V��Ń�Y�䅑��������
<�xg[,����/�B2<�s�u�1Oyx��'9ԋ���u����:���j�&M��9�'����qd��_��-�3�u��J� E�7������a���1L�ef^�������T�rh�^ch�ċ�FDXh݇w�@��6*�kO�"Ф��P�ڷCk��m
���Q�*�oe��{��>�a�_4q���%#j�PR�L���l��|�r��&E	5&�ǆ�>qޣmɟ�2ت���L�~�[����8�
��7��7X�h�o���h`x~�/��<d��0�Ȭ׃1[a���%�+�	w���KBQu����e��L^�����ȽC�[؄�P��I��(g-�2����t7K(�?���[�I3��z�_2�D���)$ӂz;H�5 z}Pߘs��C
�&ʕ)�E�e��^�	<���!����7�g���Az�޶i{����`ww s��^�_���w�����?e��dKۀ9U��gj��A8�ݠ��,��I�]�E=��z�p4[�޻�F��2	xΞ�,���?C�7��Ԭ+2`���J�}k�^�qC S@c�k��z�]|g�Sk��<eU�u��)*�N���U�Օ��>g.]H�����&@�v����}`{���	6�STK"F��4����r8Y.;�k���ZT���?��T+`�qe�, Qv���o�p�h��3�{�D��[T�ۡf�8�
�7��o�Y+�/S�aZo�$2��=S�[��ɝ��%v��,3����]��v����r�ʽ��r&[$W�{�=�>��ӧ[0��e5�)�� �w��qE�3�$����][]��<��"UJ�⬂������t��E��[�)��&j
T1�Yâ��GM�B��ԥU`L�c�+^)�7�䰇����T[���_�\V�kç6�&H�H�k��0�#G��V^�z�|N�����2��0���^S�뫷=M� ?wq+�U����B�#4���?���!�.��4��T)=�=�%��������m��h����Eе%��rSi�!m�����g���fc��� ��j�6�<�ҵ�'�:��0�L:/���cCn�l퉽�A2���N<YI�R��Jf��З�3��(���x�]mZ�s�	7�CA��b%g!�AK*P��rvݗ�M�������9\��+�;I`��)�W�m�[t��R��-�S��W�[�pYl�k#*2)��^T]���)u�r��1�m�&��2�rJY,��0���kK�QM��J~KȰ]���#�^�5��*���D�Rbŏ�Ik;%�h�_m.hr�S�b��*���'���%��l�����#�nӤ��[��I�؜�sbg�;!��"�)�)��I'�$^9��9�sSCdȤ�v��iǛv�	N�Ƚo���d>^+����coX�g��MJ�����*.����4��3���6��b��φ�I��e�����n�_i�>�rR��o/F��\s �2�d6A=�M�������=r��43�����HY���l���"X��ȓ��?����A����>L���E}���a��;h)T��Gz��.m���ay@�{+���vPq�	U�!N��(8O�[�K)h�pi��&2����`�I�v$�WYM5w>��H?d����E-�q��z�·��8)i��0q�8k�<�h8������wb�|�j{���}[o ;�5��)���qj ^/
r?��Z�?�*/�J�:Z�I� �Ӌe4۳ ?�|��r��6+���*�@�*:�2��X4a-�xQ�U�/�a2���)��р���z]���@�J9�ػ���-#�[�S���&Ś*@��ҧ�4�� ��5hJs3��y]���Y��>r�@b�yᳵ����~R[q��>?�)���{n��uBo�ՀjH{R�?r�0�p<�%��!s��5��xz�{|�˟���\��wLX'��J�65A�jضJ�T;��y�(_�A�䱈
mu��V�9��Ӽ�Km�����'`�0..ױ��0I�� ̓`3�'%�F],P��	��qlIw5���������10���tT��xe��}�÷��L59��P��G~|`A�HoT���'%�����/����oH�Ԃ&@���;@�:��ܵ������LV /�ˎ.��-����(	��=hǂ���,x���Rɭ��D3H?��ҡI$d��G堥���ckY��~Y3��^(�ш���$fEM�3脇�w��qg�v=C�
�R���m�c�Y�nvb;�V�A�x�Wx¾1���8������6� P�����Kѵ9�]Eȑ�q�g����c �*q�Ȁ� �z��s���Q_-��5�uz�kt�g�!(x���jlt�*U��KW� �_��=��;���E����m��*�-�*&U5!���,��.�� [d,��`�����x�d�)Ҿ�0������)��W~�Я�a�F���oȵ#���J.����M"odJ� e���
lx�6_�n�y�QX��fL���fTk��%uQ;jn�Tn����&�S�N9�n�=Ɩ�柹��YbM�E4>��S����V��������]F�Q�%����xǰ����cd��Y�\d��V��-�o�����1pe�E�^���$Ét�|ѪR��nq��������+�Ud��j�4w����}��i�vT�wB�{w)��Ú�f�L*ơTA"��Q�"~�����Zx�~T�Zo�g?A�S��bd�S����]�!�-e�>�⪶�=�=�R~��pQE����;�� $��d|x}��L�ϱ�c9@U��0	�MnJ��){���}9�w*5����V�t�
�Ue#�����5/�X\HKd�\�b9*�U�{辧Q�
�1�t���OG����7��h�ܕ�Bb�$�j��d
|]�g[qs��սu��'��S��������;z�j.aT�LK��Q��]�$a�k�[q'kx��æ5U�C�qԍ��m�@oe�,�V�S����P�z��l��?<�7���1�u��nC7>�Vׂ��'�;£S�#]��+Z1c�Ϡ*��Q������5����0�xe�,����ݡB~ܩ$�U�ABm���� ��CSU��Ix�y,|'!c���r�ĵ dQ:��tJ8=�F/��)�m:�%��$�_9'��A�]MH�Y������ߧC�e�	�[`D8��jda�ˀ�~�Q
$#��b��G����0Έ�l��8��:�J�@�;/��g�!�Q��J�$k�Ztm���$�-W��(Kc�5?@Z�(��̴Ү�{����,-�_tKɺ�z�l�����*����#��K�%I��*-���ZQ��O�O�˻�^� �4(�.��P�0l/����ܤ��
q���'�,�|���Ӊ�w����q���'"�D^�ph�@����X`����!������mߨ5����u/W���fx�/_m}T�Z���ְ���nğ��#�1p���D��1�bpV��Z�����pj-�g	h ;4W����^�)��v�#��b�x��}����N�o��	%�~�V�}��>"uh���r3����6$WA�m�8:��j�5��t�ݫ jJ5PT�d9�'~:�J����y�D�铙��lϤ�N��8��J:���`o� �P���	*q��H�'U��5E[��}�64��:�S��P�x������G~�2wނڮ*Gef�M�j�d_7Eϣ34֐+F���b�b�$C}4������3�D���yn;��
(�{�����L��e��{����Hg�7��)y�:�8�0m`~�B��������Z#6��Tg���-����s*�끱��<T_0�I�H9e�cL?�ttJÄ�@�ZQ&i����� [��}F�͖�@H��6e"tN8_F��<���{F�"��Bf��塏�AH�n�2���ǝ�d���{�^�ꤗ�V)�:R�ZΊ�n�t/��@�Ӎ�ѩ� �Yͅq�C�����u�']D��o�}?�më��e�?��J.m!���^*�}�L2,G"�"{��@�@�b �'��<O~V�BX�h��$.����a3����`�ʝ�͞�˲�7Z+dG�g�%�J��Y��-^�j�I�|V�1�3X�cga��A�X/�F�<�|���N�
���|��3	��.�﫣9�[�"6� �,m#�X�6�բ���2k�������^O�`�X��L`�ر#)�R=u��
]�n�m�Ś�O�MV��&{#B5�K�4�/oJ�S�}pH̰;��F1(z?%�*�%�OL���g��8OCv�a�+�[�ş�ay��lN)pIxlf#k!�h�F�<��ȡ��:�~u�w;u��%H�M�+�T��o���i��]���~ja�� �[��R��ԴO�پ��ʃMG�X�ݞ�B�g{W��@�LK��}(�$���+�4h�`�����D[�����t>�*1�܊����$����E����Mb��8GXR~�Ukd��x1�yWǳ�*�����<�/3��̥�I�>g�[Z�0�xv��*�q��nb��]�Ǔ�tkV���0#c�_�_��ifA#�9�-;��W;2���U�C���I$X�l���� ��u��/B�?Y�d��zm��F�t�l{�q�L)�����ݼ�t�ѻ�>۽O���$'�u�&l�(�g}D>��	)�L?��A\F~����0�e��t�Y��p�3�rZz�гc�����F�c��хoV�H��MɈ�N��Ԏ
�~jK��č�Φ���2��ɯ�b���`qMSH'v�����X���2��9�F\Ȫ���]6��}&}�:-')�Q�*☱}�;＝,�qNx����fp��h�f1x@Z�`>xq���3(lfE�~F�������� J�-B�!�C�^���b*@�a;�ʢ�%3�����P����x=-(ی���;uZ44;�R��S���}v�&=L�R����w���u-�";r�n������
V�Zd�'lh9�?�.��ZQ��H��l����]��%�;]�[�� ���׿&�{\����Xǽ�a׎�0Nϟ�%�o�ڱ��as�k�3/MBC}[Z�R_&F_�t��S}��mw�Wr9Au�O�D,8��P�Ǧ�Ŗ��+%���o�~�)��5iL�xiFt�6l�����%���vbL R[w�w*U�W䱠���-�ԪDM�8�2@��+�{�%1a����H�-�~�L!��v�
K�ZC�:�\���m4]<�n��ߒ��4_g�nm!��5�s_�]�\m��)���)���C���@� 1ʤ��-� g�
�,M?�Xݱ���~��j � �'=�??��4�-�B�l�����>�z2*�@��g͌ubEq�Ap�-i㊹XK���9T��8QqH:�L&q҇�Г� �����uޯ�E3p�G�0�e���|zbf����T
tj�SX9�����r���z�[���b����x������{��%R����
�|��M�\�t�����z�jE�ju)7�7�� �n��c�w�oB�{Z[u�>+��x�j��	 37̨��A#!n}�Y��Cq�rgۂ�F�ka�M�0RPuP�q�f�o3Jc;�A������0w!o�f�1�l�YE�5��A�W���f�� �0�������$O�h+j�/O�K��1�"���Ꭲ���v�S6,6����������mB������?&H	�i!�-|3��'����"+�	�~���S.}��5z���JPj�W��zN��A=K��BV3�R��.9����J���Jk|���J��kh_�*(4��}jC�悈�p�קv���&
����`d����v��n7o�Z��L�H�1ČQH�iB����}�i(my�b3�r���Vg4�fQ#���pD׆AG��5΃��>���t��(�y�[�{�۽���pk��蹩��ܣ��i��j15ak�g��`�&k���u�Z�o��ӧJ���t9�?�3b�c8R���t7�-�ԝ[ZjM(c�xl0��?/�n��FW�>��Myo$��;���2A�/�gN=Z�*O��^���5�L1���� �曟,��T΍S!�T�$��:���D��Ħ��"��7<K�ԍ�9&��`�(w)8t(xMQ�	��ƺB�k8����DF�_�S���\�HCP'�'`�SB}�8�(O=��l_���y�+����qhn�l	��X�>{�I�ڝ3.\SEP�k�u��r��u���+�r��� ��1��#���]��0����%V��L�,{`Xc�sI�z���Ԁ�o$3�Z�h���$M%�%쵮�Y5� ��&_��+:���]�ܿ��VQ8M��m�%�o�=��z��3�Q1���8=���y9�O&��۽�C�6��q��%�Ji/�e��O�g7��Aa {~i�"�6a���"?�/i;�q����IG�@��_�!�JA{Db�A�>H��W
R�!Ϟ�Aeعk����Ln�x�Q{r�a)C�{����3g���b8��#L����kI��k���40)��?K&�:x�o1;q|[޵Vϵ�Hb��)�H����Q)�p/�2N^�����IC���Q�P�u��#�$[�1[�f֜�*�Л�@�_�]◈)ɲ�]E杞	�:�>�xЊ��d�>�fB[�K3�!A��U�J6�\]�}�P���e�q5�O=����v���`�kGX�Jg�iͳ�b<	�aD	Y�@�R��'$����N��$�o��e�����6�"@Qq/:|:Yߓ��7V�y����.e�X��<;����whe���=��jT�F�'/h���":�o�k��#�z
�FIj{�*��2�mϵ��a)�e�)�YBU���/�+"�����eK�j:7��n��z���BI���0�W�����^M��X���80'�\=�A�>E�X+�,��a�Dp^v���I^�V*b[����bt@{�9Z'A��xzI���6Fl�r`�Z),�m�\Ĩ��?l�)�O�x4n��L�+��������j}���9M��/a�J�6- ��pY�i�|-�B�?,���7�`��)��9�����FU�Yq��� ڽX�9v�-]y�\҂�BnN�Vây���)��3X�����>���)�ᠿ��c�'rP�SV����!�^�C�C���p�'m�4�wI�s�7}0�#!@,.�nt�|�SE�q42�K�������n|����AiI�M_{�E�q(v���=Dy*�_�B_�#_>���~�W��kp��:�A���ٓ7�ӌ�رP�} �_b������S�/JPg^�ܜ�	��E+���`{���(�\MђB�=�r�a�Xu���ƛ/S;����H��p�/C��j#،z�
Q�G6?�ϯ��i�_a��J��$~CYC���qJ
�9}��=���d_l�/�گd�l_a��O[�
�˱VTS�[�GҶZ����٫�IO���}iɪ=.*�:����'߹a2`΍����w����I+~A�%�.��(݌�#���7>���P�9�@���2ѿ�����@�V�-ַ��l��F�_F>Vי���i�EYޚ
��H���}>3�M�P%�1�����b�*������VnG5�(�~k]%��F��`�� "y��[��{�j �
D�r{�U��U�S%(>��(����S���	s#Z�^3ll�o�=�
���E�"[>b�.�g�G��t��#o�t���̃ڨ�����s�e��ϱո8��L�%-⤳��*�v���j}�&nT��G�Oȇ�x�L�3�%#eT�BN��-,bkJ���g4�؅t$�L��>�u���^y<��bZ���JK]��vA]�Ь���h�oS� (?[�~j���*��!�m��}&)�+��w/�!^��D�g�}!�?2]�3}�4o��~ⵕ�q��ځ���&��_�����H(~ �,����λi�Y�u֠�j�n���exϚN���@l�:S�]���΋s�l��CE+����j�OK�3CI�����>���'9�����Y�hì~/��¼�D˷+p�yL������W��4�Ho�_i�L�_n�-�/�_��s���8���k��Vr���#(T�d>�[:q_�����ŭ�n?9������iu��Lׇ-��OX&X���C3b㖿�q*�cy�X?>�2�o\}H��*ģr�p�j��zTA^��V�ϗ$�)�{���|cj���|B`�n].)�w��8Z����	'���� "
F௪a:���N$�{���dǿ�@.�X�1�j���a�BEr�O�I�uk9B�R)и���5͘��C$+���#�_�<��`��Ƒǖ��-v"�	�mC+h�tm��ǲ��L�R���2{�Ҭ���sl�uhوE)a ���Li2ߪ�=\����{��{p����ȂN��.���s�"��'�;��ܚO;ŵ[i5����R+�=�:�d�CMG�S�mj��n䪴!G[͑Iz�����_�]p��&�Sqz�MO2&�x���m��m�NaH)����#�1:(	��6C�3 1N5��1�H�[�wT]a�5�BOb�\�b�/����0t�ߒ�,�
�q���J@�OE��F:�˔���t$�����<̲mV�D��VfF,�w�s����?! �������ZY�3+���4ї7,n@ت����o׎Vk���
ᣓl �A7Mq��+r�������Ĥ�&S�nΜD��'���~8�1BT?a� s��p0�r�E�wHuڭe�B�ZDur]-L;I+\����/"<�P�
����RU���ee���^]�v{h���Y��nD��j�=�ƴ��	��9JڟkMx����OC�z�hTB��ZG��Jcޢ��5�
�):5<�x)�n�\�l4��f����b�b��.�34V��UH��{�%����ŮT�5���
�1�,�\2�L�t��:|��a����=�V;x?3���A!)(t��LՏ�W��*׉�@�W��~C�ӎ3%@���@f��>F�>�df���c���S�p����R[2Ա�* ������0���_Ϝ��ZF��K�_�Q�^�Z, �reՂG<��_(�~��ؕU�$`�1?x�Ј�e��?h�'���L���-G7�����KI�}��{m,�0������;�lK�K��3	�@"TF�7)Ӥ��� � t��l�!;�:VټO���i�= ��#�f �J	Zy�̦+�VS�I�f��5�Vs,k
8:Q��D^�^<[��Ĥܗ
�����:�n�m�-����D�p�壡�7/5�p|V�G�J�����oJgp�ɺ1��ՊV�1�Sn2AV{�hn�i��L�����,�� ��{kr�&������mX|`��fP�����wqN���@�fG��`1]�hK���hP��0���:�턝��=wv���2�m
��UxB��v�%��s����Yzi^��/�<������/]
M�T��$h^e"H��)8�q�jI,W>���l���4��9�I�j�w�O�.�;�z�7�&?���2#ءU��X�e���n=Јo���C���*л{cdN1�z�6�c�}��-<�Gh>�t��yy>^o��N�T���|l"�O	KG)�ّ�֥t���ϩ�}���������H�t5�$,	.�v�x�}9�_��6����h������c%sN�(�9&�#�B3mM����!Y��L�V
��ޙU9�z�8�F�e���rj��#^=�Y��
���y�5b�߻إ�e�e�n�3ԓJ�qݲ/�1(�i�<�ۺ"��e	�㬢��xaT�>��A&�|O��{��?j�6�U�M�����DM�Y����Cc^�kt��+�+�Y�������k�7����Y㜰:��N`8�7��>�/���*K�&��$'���$G�"���\�U�4��z�O�q�kQ�7�D��sΊm�NT��s�c	��Fѽ���Z�Ȗ�����I���E��n����6@��6�}ʕ�Չ�*�ގ[����
:���L�0
R��.�	yy?�(� �����o��(��OE=�7x��+L�D���;O'ۚ�,�h�=���g���k9p�Kzm��l�9A!I�܇L�M������N���co�m;"�8������Mr�^�t��E[��8�O�/Z
�s�nʰ?��Ҁ>$�+J3L%��@�p�{ac���jRom
냏�+�/lb�@S�}�ID�ѥ��z;�YT�ч�-<hЈ�K��r��ɂ߶����a���|�6��~����x���M׋�\�ŀ�WI>�|/o�h�Cy+&���$�	��ms���{e���0�Vx�*q���kG����l%�L]JϹ@m��b��ۑ-j��A&&�z�V�{pUMD�e��R�)��&jğ�8����a���x�Z�5j� x������Ə������e�A,V��+�N�=��2.�K7���5��E=�,��u���<�D{�s=��]�R����ƃ1�9��� ��t�QU�F%rJ)�1��� ��aяȟ��x�~K���J�V�C��û�"���4�^i����Ŷ9�R�lmM�3����y嫤u�E�2�>׿l��3m�i��	�;�{U߼�,�!�w{�K"@�_1Ԍw������v+�\�e���W�Q�my�%�cߡEϸ�oލlM�����F�E^|�����
�����o!/����k�J�|TL�%K�H���Dv��������$� �K"-���r�ͬء�>��\7�˙��_bG��rTҨւ�JM�TY�Y�p��ZUf꫍.!.�,:2����B�I�1G�>�*�Kw
uiJ�W��w�< �P�U�&.
\}ޞ�8}�C�_?(�6z>��@�ƃB��b��4�Vc'^��v��"�{���R�0�o+����2
��H���TL�a���udX,r�'Y>��c�&~!J����������]MFQe"�"�֗�zB H{,�ݢ�p��$�+7;f�̫�V�ޔ�Ԝ�(��jM"��Bn��~���:g�S�X���}�|G��c��ek�o��+cyI,X���}���pG��Yɔ�]�LSt�WP�HȦ�)�����*�1�0��g�| g�KCgB��NL��w�@O��!�-#���ϣfp@��G�Z�(W�� �>��{C��U�i�$n���A�
P�g�����7�9�7d �;M�Ys��ab0mb2^�4�Y7�)��?a'�3J+-��Y��� �^�[�4������%i@G��V
G3���| %Է����LT�D�:�xmM���6��<���%V:�d;7�� un;81V�q�okz�&��:�5�[�}��Ê�0$�l]"�ŋ؉WLk��3��._~w���T[�t�Hwz���h欿kd1���-��<&�Y:�S;�EW�>v���s�.:����JFx:��<��Aٮ��Ue�A1�&˚z4����;�N%��@{w�B~4P�=��u%���:�s1���m���E�JLi�k�R�̀Z0���`�JR �^��@e�lG��Y����ud�)%�@���sF��ӱ��YC���'N�؝͈�/7d�C�+�{��N�p<��ڿbN)��_��V]3AC16vC�_��Q��"&��M�7u�mnR��{�o��{$S����U)m�D�I��} ����ں�)��M\;Nj��"*"xd.I�9�^��Y>�@W�����g�|r����q��t�_sE����d}�6m�l�����q-��G�Z�B[ύ�2Fˮ/���t,�+��}p0���gĚ�-$��a}p0N������l�
�>f_�9<�h��[� ���Á���}�0:�!ǰzi%��V:8�G���T˴w�S�G҅}J���Bp�|V��W��=5/eÂ��vQ��p`�D� tTS�8������1��sG�C�}q/��?��ݿ(�{�\.�sa����5y[�t1{�� ,Lk��G���&���F�-5��E�B���
�>=�
T�؁�o�&����r�����%M�-����LB��S,�j�XP��]��L{�QK�֧/��_m�;	z�
��޻�~9":�l�)=���Q�jmঌ�qd�Z3���xCg�@&��=9>�e�i7�2�/���jN!wS(ۘ��%�|N:b?��G�p�s�<�as�/�����8@��8�e�PĴ��jXE���F�*|�w�,��M��j�K�{�
[��W�:�=�����K<���#�i��n�rK��eU$C/a�{�a>l�����
/N�Y�jU���hM+wa؛�q��6H��t�;	?�;�,�R�π�Ɓ������*7�h��y�Y�θ?������YZ��p�
ϦP�}�����K��r�Z)���yߗ��+���	��~��Zj��+k2� v��~K�F���?��[�0*G��>(�7���<�C��{�!k�:��	���i?"��f>T��M��vg�F���[��O�{���i)�=�\�m��B�d��l$h�M:��~�&��̣���9���}OۢfW��ChY�N�34b�� e��e�ye\DOj�\���Rr�cX�G������?���e�%\D[@�"+i#��vSк���Z�;�?�X\�T��CD�%��Z��@T�v�VWH��Z�~	�0���#��P$�k�Q]m��}�a�g-�=��nX�o�}�Eo����r$m��<Ļ���ơ�r�T��Z��3�i�o���6��M����B��>r&x�3_����ioF`zÄB>j�'��H��\P�"�-љ�v&&[�G��=�kM�ʏ^��u����Xb����d��'[l+3���c���C���%#(��uB99���l�!Vܦ#5ʾ%ȹ%Vo=s��;Vd�#���o�%�4�[$u)�w�'��yuʓG��c��R���Rw��l dT����S�������ku��3,Cҭ�8e��ٙ�c�Ԩ�܌\��)6��ɵ~�)���+~TH��w���;�k乶CvXf���l85ȹ��}�wk���k����è�Q�8�o�!� y�d�Х�	������i�:���n�S'����Z��tT��W��f�a��*%\�syd��b����|ty|�[�c�}h��I?O�3{v�x�P�^�dDW{���!��_�Y��ʣUL�ף�*V͔�U�(@�*�_$B����1�������焵��2���-	�ArA���h����������R�M���=:~NE}H�_c������wi�|n!��^����&O�g��1
��?Y;NA�_0�����%ϟ����j�DE�яh�3�ˮԌ*�}���k,�͗��fmN����s��T7L�@ۅ��4��W���+�p����� :3'L�������=&���p�7#��1��blH������Ǻ�����/�b5�\�R�9�_-��.���n��`<�J�`���\�������V�,@�q 1Hrc.��CLddG��8g��6Q��F��f���5. �����?Z�f1)����҅+� �1h�VR��Ţ��C%m'�ܘ��"��kAcNę=��96َ:<���o�����~�h�P�`�J�Ք=j�PӨ��P�R#��D\aQe_$�Mq4�]a��l9܁M9Z�ĵ(���Q LYF��)���U����2��5���$�w�8���2K���a�@�E�t2�
8�ٚ�RW]4��Ò���Cy����ű�����V���Z�ʯ2C��f�#7Mh�6g{Y�d����ri��ԀśW\��fp^�7�Y�j�g���O�9q�!��7JZ�
Ѫ"�d�@?J���H�El�˙�T1�;R=�(_u�d���XNd����s�:��q_<�0���� [��޹Y^*iN%�Zm�D�B�*�(7贮Ңk'�KR����hp��қ8�s�:1�[1�y����c �����f'���iF�-��N��3��98�B��1�mL2�6�
��E�?���'����<��l���:WHj9��V� 0���ӳ���Gf\_c� ��T��S>��[��4VB?�b��j�Ğ�4I���8kM'Fm�fk�����(.¨'ߢ?�mK��Qsn�#��*gs���)�e���5l�I��\�|��9>U�/�0J����Ӌ��X�pLBs��K�0<�G �d(N?�^�_���n�6���J<�K�ʞ��f��3��� ��ƭG��o�|�Se,��&�cdAl5�!���mu`�hA��e��D3:HzO�:,H�A��ԛe�"�R�8�=<���c�^럫Ւ3�����U9�`Ls6�.�<̊�D@t��͚�eaT3[�k���;��1VCd�ξi��#&�O�xկWh%��]�����Ҡ�b9(O&#pBN�cM}uG}&8�_�D�䳩���Ȭ����f��̃PޫJ̔�΃�Rg��4'���|�2�(I{0o�������x�ZoMkF#�x)� +�0`�ٷ��.1�B�y��}��kO05fh9��Gp�q2gp�W�esNʄ��$o= �H��*�)��[��W�l�õH�D��Z��I�Qg�j���� LO�q���u�Y&�j�����</ �_�IM���Ϙ�]
�a��M2�2��"j�}�j� u�AR��O���x�D ����R�=Q �Њ����t~�f��H��� C�������
`��vPQ2W��ݓ}L7R5��,=����$I�a����*Cp����L���8��PP�+!����/,/�����#���{D_��2ҍ$�2�}�̠�k;]P.�((/������ �(������F[�t�5����9��&���bh���ۣ�����s����W��<�E�啚j}-�1lu��l(�\@3���ݴ���:>�*�e[���u�م��Ǻ��^8=w&�[+��������[eg��X	 i�D����k�����g�+�MR0*�Y|��4x$��M�n𹥝�7(�ˬ�&� �Å7	������� 4��-���s�77|}�ϧKt�n���
b~��E�,�_�'��l:E����jQ�]�n~	�}�lO_x4[�1��L��x�RT�p�h���J�ל���	�d�Ⱦ�V�KA}���;�b%����r���P6M�30r7<>��$��i���0��@�(���?Cj�p5]���&��	��3(SZA�D���u�d���Q�9
\�LU�Z~�ƻ�=��L����`ڶ%1q�6=͡�5@�>ύ�o��_�%>_ֳכ�hM��r���P"�Ě�#ɒ<~�����Ph����G�뎺xh��C�����"� x�
�zb{���I�瑩[a&rmT�S�;1�����]��'8+I��+E��Z�B��Șy����2N��&
|\̕P���c9���o������<ף0��GB	̆"ڣ�����T�O�ڏ�����L�����67cW˒g4㥅�I�j�~�x�*r��^f���>'�vQ)�nO�����J��H��s�g�0�i�� uF�r�9b.�38���PJ�br�5,�*h�wq�#.�d�u��)��V��������*930-��[(����%��l�yEk�b�Gd��
�1l/.z�~�a���H��'2Ƨ֚*�l��2],Z�~�?ഭ�7�R���<l��U �m�l�L�F0��-6��?Ľ�G~��x���8��F��f^�����5  �-��#D�R�Xش�t^��=��$cȐʥ	���J1��_��5Y�9��� %L�K�/�!�a��B<g��}��M�+g|}b��"��;��9��I�X�����W���1�w�h��P�a�&[D��9q|�s6S8/��8T�`�!�������˦;D"�˨��Rb��R�^ҙ�O�g�� (�\2X:��Վ��Rj$�Z�i� �+�̲_�|�����%_���$�4��0�(.����hrs	}R�E��cc��"�v��a���� ��!�z_�QI�_a��}}� y�b��-��C��>��y�6��,��É��<jՇdE��� vD�߮i�F�B
����B! �T���8�!!>��0�Ǝ_gű�T������)��7I����4LaH��v�E��Y?�cM҃�3q1�F{	X}2���Ѱ$n�"�,҇�-����T�a=��r��8۱���G�_��1�#�ts�\�q%nk����. ��2�
�^:�\���MR�����B�y�BBO5{�+��6��Dj˿Y}�9�$j��돜��h+�����>��.X��^�����'U�r���nҩû��sZ���H\��Cs��j�r�)ҏ��':}�C:ξT:lf�K�T����Pg94��;o��C��4������+�-�/<�$+).6�~Π�\�|g��#��5�0��&@R���<�ne
L0Y�kW�X�D�Pଆ�g���m9Ō�>f{4em����+l2���bH���5%��Q��D�OT�1P��گ��%�ʚ�u�T?˨���j4��TG��6�?��^��Ø�}�����ɍI��'c=d|���H�<��Zz4��F������΁��,�΅ް$F?��q�{-�f=����� &5��W��x�NJ���0���z�b��n§(�wW�������a��Dn4�〈�{J�������jCDg��������zO�&4�����/��儐�L�{NB�����Z�/���%�e�F�O�E�%���5XMO���y+���P�w~����n �we���ֹ��B��=�� �D�9`Ʉa\��2�:�R��~T�`�$�KZ_�6|�op»6�%��7���m~F�`R?EnVf��l���b��ĿR;���Ƚ��o\�ߴ����U�ӏ������4����-uDs�T�U(xK��x'�ѓ��h��EEO�,��X���/���{��/P�b���^����jF���q�A�Q�ַ�>��jv��g���0e�;���Ҟ;�>~#P��w;��
�sB��#fQ�ҳ<G�n?S��r�*��8+�,Q;� ���E��+-��݊��-c>�{��703�Y��c�<�����j�-	1�L�8���l��t:�^D	��OK+F�v�Ji~�#�+�ɟ=���{ϳ�'�{��	��#3��>؏N@v>��֭)�@�sn�tl �ƕ�rv��\�t�d֛���&��|�+����=LT21��e�獥�]�C���ZG���Lť~���1�"Gz����1Q�J�}���ƌg�0����Oi^��l���6@�C��
�M�o�0�m�#U��-����������#ڙ���4�:A�>>��!/?@%��>N��D�.�A:|G�)��Y�c�����{�7�6P�%Qr�e�u� K,�D*� �zÐ�>N��Ԗ��n �%�D{΢μb��� h�V��*�	�f_�yo��$�0뽵"
�A��>��L�o��:>+�U�RQIvJ�=ެd���4��1�\ILh:��mr�ݨF!��Z����GxVxl�T���ņ[s.����K��>�yYl��{bH	U�b�Q_w���@D��z*��E��FƉW��Su�J-�"���]i�$P�K��'��1'	Y�0O	"v��r=D��F�u`j�!WL�^+X�=-l�^��)�T�NE�jm[��'tH��S����R+���H������0��%��������I�?����9�3�[чyNSj3ȄO_g���w�u�2�\��2����%MZZ�"����Vۗ���Sv dx�ӫ�WLUr�Ik`��Eɖ���Ń���1uN[�U�)���@Q�!���:���E$�8�[M.����\���IV%c��6'�n�Z�ʄ}�ŝ�R�ʌ@�Q1"���x�v�`�a�����ִ������o��w|7�S;0������0���?f�ajk��3Y���M���Y�F�/�;3����,�d��u�����e����iR��L���5/�����8�V�I��М���-�yPa�餒�B�O�=��������� ��|��n��	�M���^����Ǵ%Q�[���@��h�h�^`O#�����[�����KI(�_�k\+�� 6�}sL�?���o1�7�b�L�2by�H}�1p4��iR":A8�R��I ZR��T��P��üR��(��Y�����S�+k|B��2��kb�p��b�q��Bq���ԫRͣ�Wld����<̻ӼJ���²��Y�N�/��lv��^!!����`5�k���_ӥ�'$M	F[^r��Մ�>��,IݢG�h	D�&���lqS��a�X�5�s7��K�ޚh���N�߆��g�:��|��dn3"���3Mek�[���6�Y�Q�aq\mtCE� ��cط�$��w�J9�f
#1��E�YB���|IҍF�?�rK>�4�O�
��A~n9��c=�*��[t�!K�ErM&��$P���"����9�B��X����Ac�`5�%�>��JFD�G���Rq�]�>k��U�k��a��?I�{Y��WR���E���E)��@3��)�T����6�AF��	�~�ڂ'�3�i��b�j��MK�2�we���8H: q͏�Bջ�Ŏ������eg����j��*�:�H�C����N�E��	g�?X�B���7ӢIf�w���,d��a�^������B�x��c�9k�a��o����sS"p!�"ʢ;�1�����f�%E�1��6��	��9�trY9�\�``	���ķ5�b�g�������ʿ������͖����[wrUg=����̼��J$.vY�9~��9��dB�6#�!���*�v�]���l`�s0A�)��B1�����Vf/\�5#�48>��':t� *�����̆���n�
5���E�N�'��H� q��O���n2cBf�`b�w������ީl����~dj�8�ꚷ�n��~C_�aA�x�8�+ؖ:�(�~���ܣ�bh�G��9!m���#/!RЀe|������60��mv^��(:�hP�!�n�R�����/0Z���L5A�Fф��Vƛp�`���\�V�Z+|�ew��bm��׵��Z֞�C�U�2)7��U�ګ���R[!���Ν;�R�t�v�h���,��\��4r`$_O����O^���ː�)]���Q����粵[�`5�G���1Zo9���޶��&;ٗw꿫�E�]�O��הݾ�
;h�[^��X��~!�@`:Ƚ؛ 6��{��V��~��d��Q�"u������ZPn�jX��)Q~ƍ�k���G\']�T�,���'��d�_����'�#B�<��5���mDQ��z�Wב	��3H~ܗ�%D�рR��v���K�_l$��������,0��-�c�7 �9'!�� ���⌈X��c��?u���3�l���1�$���S��޲g�*=L�p�pt�&@��n;\�v��hi��B�$��9��\����&��6�I�+w"��_�ʻ�g�h�j@��4��Ꜹ��0������c4ä�KY��IZԛ��{��Va޾f�H��K����.�ֲ������ P#���@�ذ,��iE�c)��/�]�_���É�p�̄��;��)��(�:Y��O3Bx�s�*ɞ�e�d�ږz�.��<���K��v�[wZI�a��(�� �5�D��J��.2��OfIBG�:��62�c��-�����'ax��9QBb~�7]���>��A#*�k,�bE.n>��i+�G�ūEM�� �xf@��k�:+@���jn
��z(fo�v<��AEPt���
>�ӖZ�)�)�%M�Ii&��R�fՔ��.�Vk.W.R�/_�wQ��v�f#,��^V&���F��O�r�e����g��R�=������H�aqȚ,՘Қ>��_�=��P�Ȟ^����Ԭ���`����6�n=�E9�tY@���nM����5�z�ԩ����>mY��=�x)�	�?�|Q�}�W�b����J˴s��諟��������ߗ�Y=����vU, ��4����"�(T���l��kYԿ�g@�٦�
g�t�
0ςy|}R#�%D)t�"���b�FX���?�Um~�{$��y�M�����R�]�C8��	2y�L�,{��q.�v:�eU���a
�5���A|�C ���F�J���v+5`\ �X�~���+Yf��{��(���5TF���-�
$�LϺ9�
�,+��sR�'�958��.��VIj�O�.����W�r9 HO}#����tz����ǲ�O�6�b�[C�����\W�57f�H�T��Q�9D��b�l�z	'u���J�5ߴw��bp�IZ��k~d�G���*ZQ]�b,��%��ː|����|wr�F����5D�&Ͻ�v�N�~��:���:�(a��{9c�i��� *���� ��4`;�����+���ڝq�E�N���X끰'��)��iW��7D�Ǒ9}2�w{T&i�J���`0�oR*��������;�����kI�������)'���1����u��ڻ�N�Ȑ��S0mɎ�TDp�U�mj�����f?�|_���?AUɀ��ʭ$uL,�9�4��2����8Xrَ��o����!Y���E��j�ƀ�,��:�9�b!M�?A�`����2�`�OH�*���>x��:���oeu��m��x	+Vl�"x�����o���`UQ0
a��Е�ft	���T�5���O-�:�7���!k�B��?��;�5��a9��i����T�!�<�����=�6���+?X��p
l�"y��Fa�S����������h?��ņ�-�]��#�������M�Ej1Ҩ���O� ���$��Q�~k:#v��u���H"���gC�e�����b���*d�ф�)�cV5-�$~M�T��^ā��5�F����@���r��d��l��VU�#V7ng�5j2���Ҹ�5�:C{l� � ��xLl⽶�5���w��$�����I�}v�~���P��eag`dz�x�����NgA#S��p�s������="{5�
����ٵ8FG�Q������wP�%������Ki=��LL��cg�>�a�������K����)|�Gյ��~�^P�_�S�tz��!1�@Dq�Ӈ�a����i���?'=�e��:����>��d��c�]�JWTAn��������Y���A��ꔌ�
�!vtd�� jN7ԭ$7�G�zm�(�J��p3�q��� �2�Fk�wtܟ�O�;����_���;/
;����P�5k�֜�����G*�,�lr��[��7q"�Ǽ8�ZsPO@��]NF�[͉�PZ�n��#/���n]+�e�8F��u�>S���R� ���D�޿w�+��u�����_�|�������vd�0�á+}���RZ�?X��g�a-����e�1�.u���iT������#�[	��|��q�tǓ>���҆��s�u�V�����{XJ{X'�ѹ@�34�:e1�X�4��L>(W�l�9T.I^ux�աۄ�]�D��gwb���ڼ�l��w�}/v�h���>�e|����>O$��(�y���.1�L�}'h��4޺�:U�Gpev*�_l�U����fX�-4��.:	�����}n鲰���A��|�dB����s����>Gʔ��»e���Q�q�����/�݆q���� �	��H���Z��?Yί#7/��	����gV��� �e赨��T��:I�7k���'�M�#�)1�{z�H���0��_.?/ �G5��#��P���j���0�n�9����D��<�6��F"r�fM1����lzD~z�ȫ�M"P"~O�����.����e��n�>��L�x+��
��h��B]]0g�5�"��ENR���N؃΅�l_(���ѕDސD9*1d����7'G�-�A��g>sĲm4���w,+�,��R��H�#��Fo�vEGkik�r~��?0Ҥh�	�Wn���dF�5�i�W���|>��U�Gz����&L|N��[�;��D5݄�|��q95[x�Һ�*�����J9�2g���/\p~�EZ�x�ՁHIF��	+���\{��⿜
�d��js�v�� th<`@*�"5^v���O�˄�s^k"�O����X��cj�`�!Yd��0X�A�Uc��~4 �e�ɟ� ��� �H+�e�"~�@�D��sS�Tl�S���q>_�JRe��Y2��o{F��B�������0��HY*��#Ҷ�Þ����g��u�v6��^¨��F�3��ʝ�Ġ��=�j���9�شyXM���Ҝ��a�q�t�Iܡ�%�Ť��j��Rӽ[�����_7+O@4�%;��H+�F��^4�			܆�ئ����$G~9��`�џ��R��@r�E
����9�e����5�jA����������H�F�A�����f����*���[�R���}bR��ui�\nw��v�R� �j}���͂WI�PQLEHː��tb�$��Y���O���M�f_[��\��X��S�1�(HDmA�[�Nnw��B��jƐ͞$sT��-���e�: 6�6w�-[A)9�(��H܍*�����_�g	��B�ɔ�I��[�<�aU��㝣��m%��e����n���^�#̼��Ɵ�$iya��a5�Mg��WZ�P�V����v�#��֟8Q���d���	F�<���U�
�ɖ�GJ�1H�*	����rhɴ=���ΰ6 ��a)�WFs�5/q�"n��6���2 |#��0�$!�،��])�P�� ���D�`���2���yp�8P������&N]�Z|�wx>y)L���hL��'��-�j��E�x�{|�:�{cBw|%<pb�9�@�%�)\3tY0x��)��*�=�OW�=$,B� >uo�ȕ+�_�����؄E�)����F�ʬq�B�|�&�-�����%Q�)!�$��f�fB^~X�AW11q�4�ͬ����dF�� ����آ��NN�ž�2�-��E/
lq�zrֈa� ��_\�jߋFn�v�[�R����*x�G��Ş`��s6�K@�@C�19��+�i� ��A���	��y�2���A���7{����U�ᤊ�J�6�mdOfym��x�������ҷJsDr��Ο���!T�w'����@r��kOAJH���Ϩ����Th��[�ŷ�L�JS���y��`�k�·A�u���������Ҧ�Ĵ ʜ�d ��P�/�J���y�PA�	�_�3�t2��r'���oN!�f�Cr
��:�'k����
�j�p�x��*u��@�t?	��*(q�%y���0�E��û}'/�%�ap�WIh�-+?��M��O��"���?���ZT����RKX��,a��B.);%H�
|�[ğ����H��j����Ln�&�S���ay�����.��$��˞<y�B����_�hl3qM��9@A[vi�s"��"R�Pj#F�P����{d�g9�īX(�@�7e�I/��f��/��Gf��Ph��(�txL��`,O O�DJ��X�
�0R��9��ww%����gk�ɦz�w��S�i%�!_a���<��$�(�F�f~È�7s�� d'���ފ���%"��T���Ds޸�\y�:#n͗��3���(��?3��M�4.h�n�zC��Az�����I�M|ǈ(�8B#GPU1C*ĂqA!���#�Ӽ�t���"l���(�T\���c�9���'�U�|�1��6���[��!2� ��̂����O�L�a��El彁��h��,X�6��}26�Ҽ-X9���Ou�M��>�7Z�[�D�jypy�"M��,�)���I>�.�Z +�yבֿf�����V�"��]���0���5Ko�_��M�bI᫘�3���b^�zSo5F�0�{���*��~~��_��1��sԅ��S"�b��������>TF���˒Zg���m���BU�SgP�&���Di<[�0�3���W�h� �:S�T"��q)�"��zf9/����5��ϱ:�4v*�����Ӱ��`e9YEI]�a��j�i4�����h&���Kt���mbc�W	�G�ar�,�G�8�Ђq/�j����3?�	��$��\-�f�'�ܒ8�#Y��i=��}�y	�_=
�m_�@F�����t1�D ������
�b�H'��땡v�m���%n����0a0�:�ͽ��q��q4��j0��J�Hs��E^4)=?zQ�l�xܨ��������{���5�c�ߌMohH��AF�~��g���oJ��42��\��[K��{�R(e8:�2|%K]>Lu�����~QI������]Ve��/�ԬB�"�̰��� ��d>�2����W��,Dg�w�5�~��8�?��0x�#����!m��Ҭ@'�mù� ���l3���K|}/��d�m@ᄕ�Tv	���ǩ���3�v�l)��q�Z�D^�TY��}�9C{��6�K�� ɶS�M�u���gx4Ŭ�@�o���`��88k�JTfzz�_؁}������2k���N犇�٪���P_P�Z �ۅ�A`�ަҀXѪ���qq��K��ZZ�����}�$��_�N0�87��{�.�VT6U�K��#0�R��-؛S��O�~QIi�_#��	�������ZS[�^'h��*�h�7S'ȅ&D�H@��^����l��c�� ђ�Esm�� q)�2�7�F��[#��-ψ�}��t|MB����C��7iX��	^{/�X�"�i��Cݑ��ƱO`�AD�* H	�vA/��X� wP�n�G���������Ba�1m���\���禗�P�؅�o�ȇ1��t�X��{K7�Z$��r�I��x���\��fB��������˱՘/��
k��.ۺ3��tDC@k��+���W�W�D�yV�-�Vb;�ˮ��_/޽��O�`���C���)��߲��/���%�kR����볓��ݪ��H�1)U �ރl���H!5��V��0!~X&�Q<3�ச�0������2>m�����)Fu*c������ш�3Nw���Ϟ;Wc��_R��������5���h��'��5��}���ݪT�k�֢J�Z�_�Wt`��j��6gvY����<��^9�CQ4R�S��Xry'׾�t�r
|�� @��ܺ@��"�șn�Xl'�+�D�H��`O�O����%<��{m��m�AK��Oe%X�Ao�U?�ܺ�bmch��m���_�C�8�1PE��Xr����^i<ɣD�IZi'v�=<EI���CD@��;��y�G|�M���<Xm�N�XW#����.y���]K�~�.ȓUc��}��Si�Ä���U��\{������7���4��~�;1�ƒ`��揨s�k�0C����n�X����]!v��5FmC{>01˴,���W����6�?|h�*�^v/�Ks���!b]��%Ĩ�I=��^o���z8sn�*� ��u+������h��ɶ�e9���SSeF�[^�'Khw�Э.`�Q5�� A&:�� �)
��0�;1y�3r�ťqR�yX~������@�1�w�'$�<�4��a8�T�����.���C�I�l��]��((��+ �|8�5�d�l���\����}M�S3�P� �$Y�H�����|1�K~]k���^�����di�#�̃�a���v�R1���48;-�sf�0WS# 2��o'�c�2#ۻv�|�T�$E�ܳf%:��f�_e.�G�3�S��Y���(��v����[���\�t)Cs!Z��M�[�νC�<��1@L½X�����>JW�l�M]o��j.`��n�!�>g�:�����d�W�X�E'_3P�B]�?����F�=���� ?&3�9����䵳p��b)��@�>�<eT�>.u��D�1�	�]H�Kc6���v �ֱ���}I�S�m�;���� �9�U+a� ?�Iq� ]��[����l�
- �3͡�W��m��L4�<�Z��/B"�M�'d' u���bW���8@2eX����\���bΓ��/�9e`��f� �2�9�qDM���:�ٖ"{C�Ӫ���׆A�Bi��%9���1bGq�_I�Z�2��o�_��g��G<�y%�]�k��aSX)؏�R�F�NVn����%��n�s�,�;c�l|  $� �~9®�Wr@M��W�\�y؋�P)ed��L������t�wH����C[�'DPޖM�0��*棨�~ݝΣ����tөQC�D�hJi�\�"yb.�l@�O���ØS����q��������7��G*l=���ib�t5۳�������5+rJ,j�7~!�,�g� jқP�wO���q&L{���%Ya�C�e�<�v�i��m��nX#�TEcj���>� ���S���]eN+�eÔ�LE
�ɨ�6�{��8�2d��U+����$��jT@��/?���1-��h٥�F<�p� wY~9���GJ��9"��>�C�w�~&�o�F(�V�h,"��ޗ|��ǋv��]D�~0�<8��,t\#B�e��Ԉ����6��Z��=���]`���V�h����vOΉD���'�a�_����Y�mFH��7���WQ���+�|Q
�I��%�����Q�(�;׾��d���S'NWOь{@�о��,�C��]�7d��� +5��;�)��jt���[y�p�*�^e���q�� �q���O�*sVP�K+��A��0@���&�)ğ��2�f�R�|B8y��u(��!IKE���3���μ�Z̩��;;�5ºϸN	�8^�����O�`v��M@Ll�O�{�?S�`�+�槠�j�?�S@���/D�qhy^s�:�#�D;��9��I�*m��/����
��.�0�+B��88^@u���V��$*��?(ݿP�C)ir��h/��Dt7�̐�LF�x�Z{�/`�!�\� ?Yj��P/w�K򆌥*d��gi�u톮�q��d���;����(n�Mbȭ��%K�j��xQ25�uzD��)�&n�֌,E��De�TR�� �:�NA�m��� �C�Hʼ�������5�J~҅��W�L7�{�2a<N�a<N�i}��Us�C���b`4�L�Ð�G�k��H/K��\���omQyu�CI��мݸ!I��_~r ��������p>;V��`��^\�w������^d����	`������3���pgEw������T"B�#������*�	v9[A��;I�c�<���Sn��Wpm���V A?�xd����������/�+o--�Ө{)f}iѶb�����$2�
5d8�4xHds瀰�bΘ���f��&�r9z""^����l�����#Β�1��ڎ�ZʚM��1��3s�g�ΰGoT�����g�Y�TT��˵)�����~%S�B�ɕ�%��ۧbC����ۀ72��lj��aT�H�K�$pC����MX�������C{�*�Y�"~��o����HQHAt���>�,�p�H��Ep[�y���.\���i^Ut�.�/��5�#F�/E���SG���׉��[�T�	��ٮ���q�Z��zy���.tvƸ�}�'�jh*
�E
2۶�O��V$�:|���/�7r�D����%~�����g$�s�4���c�v���P�W8���B���v�C �����~	�󜚎B�B���.9S'��aNsr�����
p/��)%r����bW!��	���}������ǒB�PˢZ�&��Vq�G�L@������	ƍ����sB$�n��V�m�2�j@�xW�|B�J��=�Ǽ|Z �=�XǛ��R�� ;}R�Ŭ��l`�6O>u�q[��T"��@)�H�t7�um}*y�bm�7{9?�K�|��m��,�l�uf;ê��>���V��ֺl���A��~�:»��Hb����y�ޗ��LE2���P��#u���Kj
��+wH��=e��hWz�K�|�Y�p���&i5$/:ƴ7�D����i�3����A�\\�YJ>��D�p>���νV��O.�R[�� �'?e�dT�����W�W��������U]�����Z'�qm�dq����B(�(���U��/me.�j�Iz��@��w�bpJ-����-�����:�i�ZV����W�_tbW\v���I3W9�E��xs�ƨT���f:X��$^B&Ils|`�������;�$-��k�����ӉY���`�:W�U�L���WV���J��;�F����s=����Y&r)��]D"к!�����)c8�1����/�M捯T�&ݕ��ڃ<���k8�񲇻�@,a��!�|��.�Z̲�=FǠB޴����8�Y4|�������N8��1S�X���4z]�������0ax�@������<zzq��@�[�W�_0g��f��*�X.�I��f�Z�&*}k�_�T�R�I�pfL�Z�j ��D'%�yS��o�=ṗ[���t���o����PP���K4klN �Q_kkZ'��+^�� �KN���XXFU)%>��N�[�퉠�tMk4�G���缑m�?�u���A&��S�~϶ʽ�I{0�oè�<��s��/��i}�����Mq6��8l��a�B��z��I$�k�~���Gϯ6�n��л����٨�>��g:�p���ԶM#a�Tk��ؘEa���Q�3�6�GAm�����ީ}�7�߭�M��M��R��r�{.�E�rd�A׹�MI�V���1q��2�JE.Up�Dj��Hڑ���t:����X�ʻ;7�nӖ�dQ�K���rn�m��TK�`M��KZ+���;�� ���D���ݗl7V���H͹�L!e?�+�$�|��@���<��o��
P�#b���һs�FN���H~�Չ!�l)�5���~�HhJj�����}����cj$��Y�g�M˶�lm��E�����d%���od�ʛ�d@᩸	�F9"H+o_hX�Xx��J���HPNf.�b-�3�K�#���˳�Hb+��P޲܎�+I��DL�����;�a�R�����¬�M� �bN�q��xC*��mB�O����'3fwD�Ა��c�~�3-S���N�^t|?�˾4l�:�Zi����"�po��[��.U/z���������|�Kv��Xu�X��k��ތEh�_��!L���>1g��^O�4*������D�fSnX��$��	���[��)���FMmn[�T�޹W��3��U28�vh�/�]%�U�
\eMUV�@�H\�&#�D2_J��aV�����F�Q�E��q��]�8�"���Ē�����븰ۖ��t:7�����3UE�?��?D�����ė��r:�Z �8��[�ˇ2ܫu��X�]Р,>"H�S[�v���~Z_l�9��˹�Z���1T����{%�V�w(�����Pȹ�Qز�ǯ`5�L��*GR���i��ֱ"�"����=�c2U{f�z�#���H �y@
K�i��搊�S���o��ED��p�8����ɿ��:�a�:��4L�q:NW���|{�y��_e��	Ӗz;�9�O]%ċT�#_�>i���ՌgoGLn�/���UXu��И[(�I�}������-Q����,$�ޥk`Y�_콬0��Q�B�\_6L_~�?b�qo^O�F�����ӈ���^2�W5	K�'5�h2C[O]��T/��$��S�M}!��LE>���t푧.V�8z��H��&��}�z�������h�f�]0Ȟ*U���v���T��n0��.�d�QAM?���9z�}5��Vjyv�����р+ ���
���5��π4�3]����[�1@�_���)�	��W¶�<,,]�Z��hq��̤T��r����V*dT~K�
d�*���!L�]� ���Z�����&�=y%�����s��D5E�q8�	ޥ��i]�ڏK.gB�3tD~x�;A�ț����cb:�ܦ�ܒ �l�'!�zW��|�Z,b�<c�+�_�"F/o���������di����j�Itf�m�q�Z}U%/'��C��h��J�`�:���L�n����P���!f�X��nH����C-`\q����+݌ux�R�ʃR��@hϼ:�2����r8��ӂ��h�zD���'��kd�̼.GZ	�l�\sN�y*�k�=�z�W3�E<h��wF�8A���v���P�?o�	��g*h²8)9r�j
4����mF
����j�L�����F����29`p�s�ȳo3ٰ���ɓ�d$bT�hӧ�I��<�n2��]ة�����|#��n,����v��~N�'qw+
���u�����|f�g	�;b��bM��k|��T?[����/y�!�BƦ+=R�5�}�ޫ5�x�إ���3CN���;���������:�l�W��@t.�˱��gw�B;���y&�վ�嫿l{�ٕιy.F�@��%��M{�L��v����jq' ]�[�����Q�<���Jױ��Y�ϼ�O�F��O����."�F��_#�Y�����&e������J�t��&n�1�ʻa���&�v��)jI��5R����nI�`�^~\M��0�CnV�	%I�mR<����W������9�����z������|�F�*e�!�	��X=��m!؉s:#XM�u�SZ���"݀�ı����w�H���k����Y:���of�/��FJ���
�\:I�IxB������x ĝ]�U7M��t�5�m>܆�p��'�>{!��/�-6	���`[����o��f\�?��~G�˜ K���
Ch��(?]�;���P�d��6�1�eo��!X�����p��x��x��/L��Bwə3?��6�k��mil�~k9.<�ĳ�D�ʸ��-ܲ�q�U'���iBێͮ.���p&�:�Vw�܏!(
c[^�a2+pr��(�ir}�>r"��2�ퟒ̪6B��S�k9t�Rw%�gj?,���=5#�,�w�ƑNzv8�V�����+D�i��0Ex'o��v^Z�L���ew����9�o��	�Fs
��`��<��k2Ut�KY�ٲۜ�G���!��v�����m[$h��s�icT������8�p��3	���b�{ޫ��Zl	F���xdИ傂��]�V^<�O8d}�3k)�������	-��GI�%GrM}�5���{�"Mn��.o0y����>�|�zzӲ�s�}���R�=(1
�$�rCE��	���&1Z��g��W9�������p���ʳ	Q�k~ �_�[��ծ��2�d���=v�]�)��Q�v0��VcǷ�	n��Z�9�mzA���=X�@]��zi	dVZo���F�	�?���Ե6����mށ������~�?��R�MHd��U�&#k�_I����s���ed\�����M/�S߁ЪQ��g�b���F73��P��T��-�O�|����0\�G�];E����x[tRׅ#V$\R��EM�)^�����!+�\۶���{�"�=d�K:)L����Ño&�s�fs���)�|�F�=�[®u[u&
2[�3�n �0e���^�<��='���Wb�Βgz�_���� H\�0%]��P��|rmԝ��N�GϽ����S�i�F�|u�<�Ĝl.cG�`)�x����&�m�]�I̿�-�L��A����o�#+�-�>�rʳn��Q��!(�3Ư�n>���kJU!]���K:Gq����y���U�8�p���id�x��3R��Z�+,ᛰe���F��i��'(#�PH_��ɂ9F�tQIs�U�FP� �K��\3@�y��*ܢ��g&Py��j��~���4:	B���(�ؐq���[3������]9��t2&+>{��y����7����*�E�D�� t��O�T��\��2ח*�ܡ߼8�s L�&��Tu�l�L���	,a6���>�P6�����!��[�]��bc�y=���݉��H�E%
��
0���%h��~�� 6��]���'0�)I�C��~��qȃ��{�>یb���;Sn=�JHg!ڠr ����\��vo�chդZv���̎_Ym�(�M|�8�̔�Թ?�͌��<t��7����@*��s^Ur��G̾Ը�J�|�5����?���]�&Hr@���;��Bs�$]�bI?%���XJ6�`p��@p�r=0
����"�גk֯;�l7S�$f�ƷK,�֎��d	��%��\���L$Sա���������f���/1��M��s�kִ ��s�wԕ�����e:;�������?��?~7�w�\��u�5�����vVR�-C�WO�( t�τ�m�!)H׬��Z=���Ü���I���t9׎a����P���-Xk�N)8��$�-4��S�
jm��pK�;�h��((��4?�1o�GLk�p����65��C"W��{k|�c�nK��X,�ߏb�y��A���)�p@��p[���M�ĕٵ�9!�R���)�;�|�u[X� ����D�3��ˊ�pm_�iF)B�L�c��t��������m��4�F?RvK�j�M~NW�;�K�i`�uⷮ���|��H�&<Q1���'��{Ah2x�n&şK�]�g
�{�S�)�Y��b�¸+Y~Q���:4��T�.K�u���ylp��{�����D��&:V��|�W7#��:3_'�?���a .�������oEE��2ᶍ1.�<$�HM�l%F�����eB�lf܋ݦ�B�9���za�`E��ǝ.��?�j@�/���P��o�Q�퍂���OJ���CZ���<�n�R�:�w�� t?�W!�ʥ��8�>�H�I㔑�}�7v0y�kq��Q���x���(/aP�U�nP�q#(��G�$���J�AbE���	��V'�z�v�L�H�I�oA�z &F��Nw�����(2׍��$�ô6
g�˺��\Twe3��-�Cxp9UUL�i�נ7#���ʧ�xz{c�~t��Z�Y,��F`�	�K�AtObJ޿�m�(ѷ=O��0r�7�Z?�{��ӪpU��W��f��e�U�8�":�y�tf��1���+���q�:����Y=י�����\P�z�#/��O��p��n͆DD7VsRA  ��c�(�pc�F��#= ��-/o�%q�ei�,W��ѣ|��Zlo-�j-��Sε�U������4E�fּ'xf��#�qt�(��[��K�-���?17-�N�M�AO>6��kh��DON��@�F��:u:�$t,.�����9�����ݻ�h�J
Â#0S�J����}�n�M�s��Y���ű2Z�ts��Պs���6}�E��Z���o��aq(���K��Ӑ�������������Vƫ�Q��i���hZw�A�E��Q��J_�P!~� �,� L��K�E�-i���U�<�&�aV_��5	�#I,���;d��$f@d� �'R�■"�� ��ު�}Цm0�_k��쿴���pW���NBѹ^��e݆j�,.|l;[�����#$1L�A����k㑷 �4��{��8.�f5e$���yi�Jg�^���ά�Ң����Cy�Z��0s
~�~fJ�V������E��Dk�&�u��zǷ��/&0o���q2����<�*GhR9'b��b��� 3\\� �"�R̈́<Z�}���)���pc����k�h�?��/&T��.�W/�Ӏ��F��)�R�xC]��拥����tF��x��dK�����%�^�&>qH�ZB|��9������I�y��hC:l�;̨:Vm[_s��~6s�dLqY�)�3���PN�==)⠳&�W�v��s������Z�6�!��B �!��T���t*C���:�.
��O׉>~����,H/Oo�7��'q�'�v��������E����%�TiHյ'4ig�X����c��nu�Z]NS��ČI����y�'p�@*��"�wj���lwE��09tiH�\cDV����7>�숸tV��ɘ<v�����Z���pƴ��,�oV�8(c! d���J��dLj���	�$E4�bE�>Z|���_�q��m(K���;b�˲��^�2{�$�	�W �p���A�8K�JNX�mTܵ˂V��
��W�H�t���
� wP��ts�������?�]��n]�W{��]�o�q�t��y]�X��A���3u0�;vK s�l*4�V�VJ��5�tf:���7唺ֲ����҅���d�]^Yy?��4Κ�c�G�,�F35�&H4��A��_���/��H�T,�tft�rc�џ��`�:���/�1�v�ɬ�f���*=����H�W�%�=	W����%4pވllA$�H3�y�������m�=�{k�b�kc�Ed�\0ȃ]�\�A% u|E�I_#��%p����p�xnǦ�~Tݚ��~<�$Y'��i�v�M�S��5�8ZѪ]I�_�)��uP�=�����nS���G��-,L���2��C��4�++s�����5�AQ��4P� ?�� ���0�&n�v�����Z]_g#��VL�M���7F��s�}�6���U*�{��pY=P7!\��5����b��\_���p��a�~�X��j&�0���:)��Hl�cS������!E��#Y���ӥ�vE��K"�ʞ���Uhv��1Q��@u���M�K��"��ܯAj�<8� 椊ۈbА�!ΘE��Pd"7�������5H�1��?��y�)z1��E/�ӥ��S�gTGS���3�c��V2b6t�¤ 5��=��7|i�đ��E��T�H��f�fȱW��"N�ŋ&�d�� ��|9}\���y]~N0��boSR%d:��KkU�=R�f��iZv(�֬|^^�'83���rp�jW����\�z|-�k��9X�dL$`��ks��)�y-�#���*ْ&C����J[��yiP���{���,��3o��5�(^�c��&�� ,L�8p����{nL+�����h����q5�V_*�~.;��xmk>�&7D�]*�赕�NB�����kК.�nJ��.z:���A�aO$/A�/�DQI��V�T�z�X< ��C�0xs��UH���C��-� �z�~?d�l�L�FC����D��>�5*C��>��1h������E�Y�q�g���E��r�����P6i�f]w�[�:�<��o:�i�TB�`��B�ݿ��9��n0�p��-�?4N)�J�BZbӣ�?��I%�����D�W�Wu���~���CM -{��6Ր����ָ1�C�z%����"g�%81K
��\��l�T�=]�9qV��=���:�%��u��Jv�I��� ɀsQ�8͎�C��~|��6�!��7�.d�xS:�Pc����ܑ}�<fU�У�*��\��n��$�&���ݶ���*K&�k������j���<�9���I�V'�Y�m~�qT�\27�<��[�&fj�r��oѐ8L.B�[$>�n98�_�@��嫡6T>�|��:����� ٮ�f!���86������{k=�|�\�����neKK*��tA,fh"�@V>�lnh� T��|��+�&�ͿBz�͹kR*OP�i���hZ��k��.�
ZAc}K�{7^���9bZZ?��ԬV�����w�nƆ6/f˫XKN�I�@)���*�:���Y����a�R�j��io��xT����V�����m��"Ү�P^D�"Z��(d�SK|����C�M�
������C�c�E�7�P������?�[��j��W��
%&�>Y�+ڸx��W�E#��9д���h��D�q�Ѕ�3�Z7��!��]c@�.�f��dB�T�O	�klN�� L�k��m�E����1�f��`�\�0�3.W	R����I�%
A�7�Su�;�j0z�g�E�
ko>��ө/�)u*7��sm��(p�N�^v [�5�|5�m�!���vb�E�����N�#A�'>SΜ*���d3Q��n����*��[�R���}"O�-|�D��庂��9�Y����+Q�@!,����H��ܑq�Ds}��9�lV��o��M�VP/цz{�p+b9�D���ƀ0�j�5���iOEN������Z�����~]Y�oU?5�#�_�t�*�ᣟ�������.��j��t4oߤ^ĉC(H����UG%��I�� ~Cu:��}*n��=4N�����W��W�k@�2 �L䄫���N�{�/��mj(d=��;>\0�kܸ21;��V����k������ë~�%z?D����y�5�Q,x�=�W�|�Y�,-�0����"+��Mg�K��қ���U�.�p��Fo[�U�����E�-`�g���.Bm�	�@����Q��}lg6B(�8{���W�lzBoRL:.��:f�$�C�M���J�ܣ�z2*[R�(�I����1P�]��B������e��]�L�R��xr��C�J>z�c2��,C5o�!f��T ?7ϳ�s�C<�ɇ$"g�# �aF��fXG�M&Z�b�S*y,�k�tI�*��סb��68�L(N*����{v�t�.���Ggʋ�e�1����!A�0�wl]�a�&y�G��<X�ߢ{��b|Ӈ�;I����>�R<[1�~��s�ƬZ7������6�
�e}��:�����E��o��	jɄ�G����aj(���E^���/��7^>Boi�W9�#��HƘ`�2U_�D`���QUN
���,�v�yhJ��.�p<T������v�E*�Ydi,���[|Z޽���PhI>Xkj�{�����x�������a�o=M.��$3M�z9Mͦ��x����b�gȖ��ZҐLf�t���21ʸ�{>����
h"G�8� 	|��@so�^`��P��������k�����l�����������{�r�@��p��xil�%�b��LY�C�i�+� C���e75��܂1b��xt3�	Q�9|�7uܘ������d�zfq��e��|����{��+d��q�+�-Y5��yw�gpqB�B��}α`>���u�/���'Ɨ�rB�~�M���b��/�Aˍt��x7m�o`���BQ
���k�,��P,���%a4�]%U�f�[P:����5��I�r"K��Ðe�V��=��*W<�KR �?od��{��6�ɀ+�G}�x��.o��y���&���\*������97*"D����(M)���s˲c)��K��D�OE����M�9f}�Q�9U:Wlm(!�챐�G���0Um?U"��;��s8	ϟ����G�1�1��D�����g�fށ&�p��y		��$���V�������0V����]hP�;E��Vr���̮�0��V���K��='�~�NB���(�[Q���}�B�t���΃W��x?�jV6���{�5N�7\q43N�ǆM���zv~Gb(��j%���	�>2��p?�:u�M��2�U�9VHب��ݬlP�+�����es#�m�"9�ۖ��{�,�,�	"���y['$�[��疪���6Tl=��C��[�3׍G�?��2E2>�=�W��x�N�7ު��n����1i3�v}��ZNл��K���yh���n9ټ���8l�x�~�m�p=�|U8��l{W�!B(LI�ԣ?��>P?�'Z�/�~N�h�f@q����ՂT����̷@k�$�Dș������1n���u/��g����}U������&����S���E�{;=�8æF���>M��#T��ے��MnS֌�19|<Q�O��A)Z�.Á���u�Է?�r�(�ك2���!o5kT�;�M�ͪ�T��B�F}]�O>]���!���^~ݤ�,o�M��Z��x��O����t�Zfr(�l��0�3Z���
>I�GoO�[�#ĵ�ӛ�гp���cx]�J^��t��m�z&9�����=�LY	�_z��0�F��:�F�Tv���ĥl�3�	��ޞ�޸�+�����Ňف,)d��(�x$Ct�تA�x:��J��Y>�ȃՓ7���Dm���S��<�9�fb�}	=�[��n�u������>���֓r`�����rA��${�	k����L&Fr��վ0��f�9�t�E�ȏ-o=����\�4���9V���~`0Dt�Șik���t��&/��\����4h��TA�X�o#_�\�݄������I E�DN�C��X-B�O�j�i��|�T���v��I~�C��;�j�褶����k� �6F�1}�`��e�ف�Z:�K�y�@%�vc�������v���m��6�TB�dlIV��3�O��̀���pcP���2em�U�쵵� �ln�V�̛��p�V^BOY�p,4�r+	�q�O���Ǫ
ۄ'gR�RdRSh��kw��咳�g� ̯"�Z$B�Q�����'�1�H��%R��� =Xƣ&߬�<�tA(�������9�=�x�`3����?3�:Y�$��8r�y��ťgBX3��=*��5�u��PF�7|CXh��t�����'��6��i�<Q]̡�=�M�����ϖ�晘lֽ",0i@�k�.�J!�����Z�#��� ���l[n,9���%.1��S� �L�M���j�F�Վ��%��r�]���p&>�%'&�/H�GFԖ���0᯻�I�l�7�%�����?>��m�D`�V�Z����ZE�'����c�19@	��H��Hff����^+��l&ߟ�2�b��+{���M��b���g��0j.�]�\�pE�~�D��������n)wr������N
��H�x�Ċ��m�!�&z��]!��t���z5	����1��9I��L�v��¾`�V����KD���s��6B��Թ�xO�Do�!	�w��ۍ]_G�7ޑ_8���\]�s������D�ݮk� �A��et�᪺�;=��&�A�z� �U�}�ɞ�d�*�FS�
DY��-���'ST���*خ���5�R��	�!�/���~�ڌ��������*��y��w	��s@v�XX����RsxW��hōm3��|���{y.:��P�+{���p1� Y�"�?yk!�7�1�Ŗ�H�l@��6;�T�ol �j-lc��Nf��Y2�SC�|�G��1�dB?q씆��.�j_���ǐh��_���׀ʃ���\�˪	���া���i�Z
0��%KFUk����x�P~�A����}��s�~�yR�NΏW������__7�N�n�^�u�?�T�0VZ�9E�K�|�n��0��|�^�Ɵ<���Ҿ�E��t�@e62����*��h�"���L7L|�"-�u�G>:�y�KԔ�xt�+��
��U:����}�$��[��	�q~p�Q�aD��G�o��mlV5_9������i�b�W�Q �-�1�N���@81�e��A���-�N�� ���[�Q>�Hɒ���[���!��g($KA8�"#�y�.��H<G��4�+�C�A���O��,u'�Kd\���H������A�6�8o�{�������l�������W_���O�ј��e�:������#�����O��qݍV�qDct޶�qLT���f��Qx����i�r�B9���7�U�.�.ٻ�1�uG}d�检 "t�ѻJT�>���'p�Ԯ��ْNnT6�$h��#����-fo�Y��N�z�IHq��S��Z�k^�;�KT�̘�.�/W�Qg�izڛg�wD6��z�4s#7�6[��	Y��������כz�
��e	�ر�	��V��u:�)�صOa� 蜹57>���Ld��Qs���iQrk��ذ���I��A~a���ʻ�30�&�f�qYl���=$�s��M��>�?iN	&�6n+_U�E����P6[�q�
u  J�����i5����j����D}�����r�S_��'0�l"YxI��2MT��`G �D�+���F�;���q��ԓ� �nrL�X���4O�IX�����(��&��>;(�a
(UH!���u/.����G~<�1�P��WȚ^*����4[��z���˰��c�cq�I���,YCd(�282���n�d�4�p��k���`�u&�V������8=D��f�����-��l�h���av��̙��`�����ch ^W3�w���N[�ƫy��Ұ�@�Jɋ���[���3��<���z������Ƴ� �	�_m4�x�\��ϥ�,��{6<=�N�%8��[�G�Ŕ�q����7�W��4	���E@fBD@�r�K�b��[6�ckn�pWr�'9T ���"���~�"�i���$u�.�@�3W���r#k[~��_MF�jm0%�M������Vm�#���6)�ǙAo�k������LO�Qe
;���������P��7�:yB8��ߖl-u�jqʿs�޺5�\�9�2.A2�;�;����8<��$�WHi���=c����bR���� ��c��BـK�F��Ъs���t�q���y5'9Ϭ��� �I����c&iN�`�ĈNh
2�~���GIôX�-��}�&#ˣ����')� ���w ��*�������4eh�8��f�[�ڥ�g%)�_l��fJ3N�0��,M�.lBo���za��q�SN/�׏{,�7��,���+��H�W��� �H��B��K��I)���H,��%��	�~�mn���/�Ѹ۵#��Z�����6�'�	 O#dm	8����i�;�-���}
pLD��úUU�Sǂ�p�A��7�پ�h���+�`��g�0�\��mE�Ca"����]Rg�������jɇ!�mt��d�y����1c��wv.�]�����+�'&��J�3�8Wo���0�S��-�S�v,��Ӌۛ�ߢ�����+>�랢i����������X cY��ǜ�ȷ�9~f����>'�{��p��°~S[3ݿjd��]9�ljfy��^u�>W��<|����6���NM����c(���'Ԅ�E�y����]�H�N�UD����fI
�"ff���^����J��뤷]g���ƍ�˷��b.�l���c,�*J��:�S�wp*�w; ����3��dAg'Ϙ�Hy��C}�Dy�)+�l��;��ոI�lci]��~�IY���X�������0�����T���C٬TmlܖI�]Η��[�~t<���~ �`CTɟ%]�h�@?��X�vn�@��ڇ}-y�{�G�b/�#�tf����ESH�&���e�װCf�؜�/S4��	$z�׊�IO��j����nuq��c�˩�f�;
+��SRk b��>y�=9�~�����Bnyϭ��fi9uZY�F�S��¯G)=,e�����(�"��i��4�Z.�\_��&��8M��W��EC�C�;vb��&up�ƑB9V�L�|���b�&{,�4Ɖ�Imv�uӳV���读ݡ���x�x!�b�p���6 �3�(���ځ�$T��#S�	��6�!A�RC	v^�jc����9y��k���f ^.x�Q�֋\*�$FPZ�=��]�kq��/��\��H�.�S�f\u+�0Ѥ
����?t1���s,�[��o�N���/s�b��|�1-U�s2�Yy�d}�` ��!+

��4�I���Og�N��3�8_cV�
�u����ۍ���=8��gP��	��P�e����k����c�BDc�
6�Nd�6�ht	@����*}�֌�� �i�1?b <Ί-�e�3��}Ě�Euw����S�."a�='���1�ic4��7�������|9���F��
�a}�v�G>��V*�/6��B�%�������b�M�jxz��M[���@*߼q�+',0�k��ܚ8���'^��!wO�`�P��sGaZ�-la�������1���-L��V'�UH�4�FD;�q�aE-����%��b(�b��� bcr�.ֽN7F���,�(��f������u�eK+-OzU�2k�`K��n�Q�k��O�MJ�D'
0ZU�P��R� ^K\x�[��m5)�IR�X�<�"�X�4"Og4|Bhe�Q@S�~��"�f@��w�@�쓁�Q�)6<��4��
P�0�T�����aە����f,���6A�0A�����!yLqeH��l�BMH�F���^�L/dnR��xSd��a�5�����O�^�.��5��K/�����$/���!M�SM��8X�F�g�PBv�.��066	_t��[����p��+R��Dn��b��������"�-�S|C(;�=t��/��x�߅0����
�a���V���O�\�8WM_A�f_���O�q�hM���#�1u�"g'Wtro�3 ZOV �� �U�y�W�)�6��ŝt��?�d��88c�fԽ���㦚]o�"˒țc!���oA+�ʵQEl�=���K�5�
�ǚpך�� �^�Z���%g�"K�q�� X9-d��`�/�����3�]l0��	k��	{x��o<��/s;�n�J�	Q�p�/�#Av$