��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��<����^����֌���[��LiѰ���յrw�xi�Bx8k����괙�u�^��d�_o��Z��Ӧ!H��̌jt``1f'�8�֪��w��g���,�}G� �:�xt �m%%?/ ������y�����8{7��Ų�2]�O��R�y׻��Rd���r�8���6�0q"����t[�{���W�a��g�^��dk��� �W�j�_R�i�l>gp��UG�Bg�Mk�{!����+�z��0Ҩ�^-oka%�bOH�ObP�����0��Q�@�����[R��;�������3��[�$N�c��r7�M�>pP��I��@hV����
h�8��l�]B��X>Y�C��LcΌ����""f74�R����t�<[]ܵ[ջ`���h��nO$��Co����Gm�N�!��/.�g�"���]g�|Qg+繭~�#��G<F�%/,<4��T���[�\�1%���S�4��X�r�/2�]7��'���D�YN��&��<KW�q�.�c^�I����2�l���(};����#���y�P�b�g��Bz�*,�L�0�P��@ $�]!�� /���c�d��/9�P�����K�Q�?�O'j�v�; �&I�n�p�+��6�����L�ʄiQ�rm��pY�ss<һ�a�%�4<�4��o�u�M��;^��gęT���cfD��!���V�;2�$���rc����B�v~�C����T�����Q?c��kjI�	��c�x8��:�{0�&S��x�tm�0 �t���?���%��k��[�Bt����܆��x�SN�������^.vC�IEmZ���k��D�����-�@:���
���:��<k4���� ����mW�Ωa��/�R? hQl'�?�u:p�30�'�'"�F�?�	�F o��i���K�n��r�S�c?;�M(t�b�܁�����f��}���<�����3�$Hq�&���D��0�Tkc�I�Z�Ĝn�ݯX]J��	l_������=�<�V�_���I�y>	�;l�"Qa��~^��N��e����顉��|�1��`�~p�u8��$�pg5YEcy�������LH�t�,q>�9��ޜ
�������Es���b���(p
g�uYW�\�h���b]�:���Y�p	m��5�����85C?��~�2���A��4H����S6*mGӫ�F���h�(\��� ̛q[�{��/�.WU�H���σ�5܇��x�,i�x���p�ڊ�bLK�C��de�M>B��KN�M��`��++D�<�p#:��n�RW�g�Wh��vI|q������8�Ǉ�bY����~�7�(���euk���D�B_pu�|�$!x�t��6��r�x�vxU>J���ǚ�*���:�b�A�1�B���Il�.%vm[B>xU=
{EH_����h��>�eqC2��Rn�7��7,�b�1�4��qs���g��fSbl��[>g�v6�`<kH�K�a[�)��!��}������/-�D,�a؏�b~� ���:�x~�����ނD� �g�����ʑ��-p5���C%T���&8�=���uV��gHu�W[�C,P��b�N�*k �}[�ڦ��A���o�����+�%;�_�;��<%��x����-H`�8|�`l��¢��d�v!ݥ��	�-�R�Т/�[�^I�G�u	"0̟!�9���f:�G�ڸ8�eЕ��ߐJ�ݓ��shb�8��"�mJc�)�U?��rT�_��=���<ٷ�WDE�Ȳ��2��;j�S�?D@ƚ�eǶv�+*�k2{�����G[Â�^3��]h*��S~0|�D��w��U�,����`q����e����%�s�����X�s��h�ܣ�bLCQ���*����
EJL����h]�6 0��e~H*[�Z��P��f���Н��N0�j��P""��n�7��ۨk�=y���%\�v��d�-$�{���ӯ��u܄H�/=�w��z��4^0�)��/;G	��vٙGD�0%
)fP �����Ȧ�S��/o �:L�)cq�p��V��J��a�"����,eZ���'E@���1�K�u���:�^�ձ���NDv4����MH6J�ex#�-ɷ����1��n*7g�L4�y?�Hj�b!���2��ոd�9e�j|{���ؙ��1{�yv;��n����r�UA�$\!c;}`#��gfo>�5�/�g�X������;1��#���k�Gw��%��U�WV�-stL�P�@���C��'3���c���L�	����z�I��N����*�#>�MY/��Η�4��_&K8�b��>"�6�I��\���0BU��;%�r�:�C��0�޽pF{e�?5�*�?�y]VE�����Th�A�P�������n^x ���^x����h]��4�Z������F^�K�ZK�]�Y^�#*δ[Ef�W�,N�pfݘ�7�
�I�*?��X첃�e��nI��{�c����������/W_:c-�`��WBP�5������-+!��VJ�?�5�t�y(ᄪX5,AC�����&�Lasf����<�s��<��	N�JY�\w�	QǗ
�6Q���ښ��q�4��*�b�b�g�J����x���S/W詳�M��](x����b	$3&��S	�x<]�n�д3Юpl�-�؂a���j�pgO�`Ȗ)1���!�L�䖡�E��s.��y�������;3\���,���_<<Ά�@IF�b|jR�N~��9#�B�CR������9�S5_�=�hJ+��y�N�M!&zX|�{�|VD�ck�O�	��������;-1���gb^U>9'��Eh�'b��������p��x�6�r�2@�ڥ/��\��;K�i�E����d�:��f\�[H��U׹k� �HvޯLr6uZ$o��Cؼ��ۦTd[�<A�<G�Y�BGBR�������c����|	g����N"NH�:[0s�۠8��Ֆ��y��7����z��D��X��ǯ�]�	���&�%8�?�Կvj� ���+Ϯ�pY�=�f'2����@-�i�{8��SW�]�V�J��<D���W��j��؇M�H%����_5c��|�B,��[M���>��%$L���*NҭÖ�'�?:��͜��{T�( &�^,3\[�v����|�������:ϋ�k���Kol�,��Ov�����+8w������gW��0o�!�lهW�/�)vo5�m"$���Fh�H)>(E���;�R�]��Zl�6��у�2�b���tX�mfE�?��\M�SSO24�M�=�Sƴ�?<�E2-�I�KW����B��u����k�Ga�>�M��(�N�Ƕ��;G�,m^G
ؑk��y�	��IU!tK�d�W���Y�#(n�P��'�rH0��\0{5,`����}��[q:@-��Ǭة��e� ؓM��k��%�>�kn�-�dV�C���C����yJM0��.��z�2�qŔBO���K��J%4Giҙ���J S�
�CB٪�SMp�������I��4�'�HA��!$z/=]�0(���vUb#��Mexu2��u��I8$Q�GA&���C�`D�UBr�S2�9��.������E�8tuu	�N�8��:�QǨYweg�J���M�K�@|{ڟ�?e�怓�����|!��+����,ץ�TW�ak�5���݃�!�c���������^SL�s+�ȌI�V%�I�d�]�&�3�.�qR(	���F��y}H	]w�;)h���i}MuU��.�1�R_&j%
9b�q�0
i$|j`��L�ȡ4��1����l�⌶@�i}и��S��E�7��7yh�8̳\���ED��1���qva��WV� �������������a�����p�Yъ�#��٥ȅl�@X:/vH�x�l ��@O'&c�"n�=s�2��ΰ^ZDI�ћCU����䗏��^�4u�f~��0~��X���LJ<UFR��zB��ȏ��K�/-G!ǋ�:e^k���hQb��T��gޑ^ ,�W�@�������5Y�q�`-�|-�h��qr:��(*WG�H�i[yW������=�m3vXj9��@���~eREm3�Q�����6hIJ��U�`#3ze'�'���nG�Q-A7��  $wq��{-@���u�GW�q��Y���	��ސ�/O�:O"����rin��~�u����R��%z�'�R�m���ܷݰF_��B��@aY�mH^��B�42Ҕ4�*�G�Թy'*�&�>�W�Z��6�,E��ꑿ����g�ԉ���Z41$��-72.|j2���q6�����]@y�<�s����q�-��j`*O ����	'��M
h�ɳ#Ph��s��5_���:�o�R1tyu���8�;��7IC8)%L�B�[Q��E�#�ԮV��l�5w�mv�.K�'�ݓ��|<�z3���{���z}�'�kEod ��L�F���df���~{5z�b���Y��B�RI��N&���j��)[8�?�&I������B��.Iϊ��Vh�W^�^>�-xHm�� �L��_���Ys9�P���"�Z�3�����#�T��07���}w�ѿ�����:���|�$�����I�b�-����t
�o�x�l�T�o��&3Jx�&�%���F�Ul� ��S��}�7��&+����[�8P�16��2!�x�H���|�W��rЈT��}R"��b�-�S�R��ё��2���@�U$�ZzD2ӫ���a�=@Q�G�,4s�o7�O ��_3�/*Dq���8��5ei��A+~���TQlD������i�[B�Ni�Ӫ`�M�6��0�S~�o��/_3�ZΦһ����*|��-�/�<##��_�q�Z��9g�?f�e���1�-����m|&q0��p���nl8�lGhx�r��}6T�����km�y���8 Q.yGD�����j}��{��R�j�~.����$�z:XfA:x$q<p&#�ʧ�ů�U���,�#m�K�o���ZS� ^��;�ܸ�ؖ���V��h��|�����+�u�_m�8y�f"Vx­���N/�|^?�й`�&�N��l}�ko�iٝ$�Q��������!&��r8��/i��3!�ƭ�y�+����L�9�%6��lL����T�䂞��~��m6��m��l�/������[?�b#��i�߹���Xg����s�D� �w��&�ɾ��g6#ߨ�I�a�6L�5��՚���: �E��E)�-i������� ��i0	x1��U��|b�A�?7`�2�	̆�[�X_a��.�mOM��K�s�\ۚ�^�X�<��q��m�h*�Ŏ<v*�D��Y&���Q3H�
��k�©�A��xQȟ��z��n����z��+}�$Z+_F4�R�V��^���^!4��a��)RYM,��� n�����.���С�ʶO�=��r����Z��QG����Ӿ������b1�#Vxt���4^p6|�������	���*��ב�M��h�B���q;f��``O�~*G�ՙ��Czw�pY_H���ϛoH�JF����h��(i�)��D���H҆nl��#��<:�N����}f��O;�:�5f@0�P�P7�gL�L��p����k�gb֔�"C�9��$��9�ڤ��h���]��ை,�j��%�3NKS��⚁1��ᰞZԥ��{U��*9�/m�Ƿ�g�##\�1�i��E_�o�)�q�۹�tk�UT2XMԯW��^r�yT���(J"�et���:�A��fE�_�󻒾.ſ�=��^_3Fy�%TN,�q2��b��z�$�1XV�7��8a�fx����f٣KDU'D�0��L{d�����^M�1��t�����+0cFL��6��Gj$�KK�����[��>��q��.�.�'H��i&L~40�x|�l+�v�2̸���{��&�es�ʋ%�������c����-�m�D����r��\�-��W�e&5Lc��O~v���"��q��x�3��benFl1#��m���ÂJ��@�����߹�S:P���>�A��j6�{Q�����X�#Y���iG�2�@�j�C��l[`� ��F�����ji�S�d$��"�7.fmm��t�Ox�-���^V+��Y}���8�2msWwD遲�	n��J0y�<iu���-�5���+�M-������A�%�Vo�?4S��9E��_=��2:�����t�����$3L�Pfal�����RW���S� ��`}�6@��$����VI����~̉2��B�v(b�l1�o������� �Zf-��J�Б���E�׹��z�gO��"p���_��w8�F����z�zZ|Ow"�,�!�X��G��T��4&Z�4dޣ�]����������0�Rc�yƦ��Gԛ�Њ5ć��ں��L%f|ґ�M��exh!j�x}a�Yc]3W5��a|�*��9�bh�_��f��F�ӽ�D�Z���:�E	�l;(�Z_��{�
�R~��������k8�|Я���<#C�O����s~Jr �4{o���^����b~ϱ��_'�ےң�|ì"�G�w��%s�:#����D4����2EVg���'��#��WI��|��ۜ�Ό@�*���lpo ��3"Gbn*b��a�͒e:)��J���e�'�+�Ѻ�2�9Q�|Ɖg����cf�ڒ��n�
�:��hd�٦E�<J�RCq-��A�փE
:��Ӯ��2f�@�8�aEVA96m��r���诡���M�$���-eW�_��+�I?�!!�i��O�'� ca��}�	m�.f�v�LA�T1U�%jr:M��u{�g1������v�=�g'El�	<9k@=���?�F��]�B���u�^�Z�7�wC����ɿ�-$�Y�7j9�������K�(�j5����^�ε�i�?�P}��S��Ca��X���,��(�����9�h����,F��K���2\�����r���K�n�G�8���-^Z���$*
#�����Z5I'q�ށ>��!�|8��vqZa��3�h#1�!G04OŊ��grl����˄�|v�c����PG�9zT F�Λ����-
$Du����}����p�kpo���<9�	�h!
��u�WB?&��D�$I���Þl��fߙ'Z��|�Yp��Fx)l���v��.�,\�"{yJ���f*�\�����o޵��#���]~O�h�ںCp
�n�b�G���q��B��*�iHK*�ܴ!�|-��&���^�ŒL��<�s��B]���Y�:��{��xa�}�E0�ڝ��I�V)���h�HQ8���'D�y_^q�خ�z�55�-�|�`����z���k��i�v�����C�e��e+��d���Zl)7|ˢQ����Ǝ��D��-�2β�p��<�K�/��8[�_�:�"#.'��Rڞ�:���D2�מ���J|w�J��*�������ڃ#o�T�ѻ�B�C)������`���O�N�A+�zjz*\�iI3Ij(�+��2���S��*N�����&�b�%6��$m��4��Ò�e�~������K����J�n��s����FT/�-D'�Zb��͑��K�H%^Q��g����^��l%��R�_1�U������k�,�
,gT�B�
��ڮ�bHd��B��]��,%������p����3 �ֵr:	?�2����J	N�]�C&1���&����ơ���4�o°�ng/�P^�+��B���Qa|����TN�Z���������|��A�-�D%rd��x̽w�i7�B���]45\#kyo��	9�[~J���UELj����~_�۸���΀'{W˔�)5X��1�܀q�?��k�$����(C؞;OQ�\XQ;�UR��[YCJ���������LN���3,����i
�n
I*WL��p���c��2aEsd@���׽J�ð�P�����~ ������a�(��def�Ԓ�AVS����$@_ww'�u�D�z{��`AҞA<���y���mŷ���G�=��a.�����O��:�_�9�!�2V}�+�k�c9HB�t��Ze{Gdi�z&�B��D@slwu9x��k�����uj�s��}8�9�Cg�u,�;O�yJ�����?�ζ�N�`�12b��iD�Y��y6�T�D1�>��Bg�%��v�������uVb� 
��c�㕾6��d79��q��M��8�۵�W��^$:�5�{�,�	E�</���I"Pk�Ų��4*�c?�N��b �wD"��j{,MU�r�9�z�ȫ��c���ٙ�6j�WD;wW^�����9�-T�2K�4z��Dϳ�������B�;�:�+��,�j�ڼ�Y�ox����ǔ�mu�p��`�@������u(��Ӌ]�C=�LR�Z�ް����L8����z���M1������!o�]��Y�&	�HrH�"36�n�������
ށ���9,�(��?�g"�s�v+�E��aJ$���Ö۽������}�'t�L�<T�ғ!������E�	` ��7u!z�\ɜ���`��S�Ъ�d���� �EӉ��NȘ|�_M�L�D�U���"�	�/:^Ǆ�0N�;�=�<h��� ��ZQ$�zSƙk�XOZ�G��xE8�2��ɠ▟�f�WJ����w�k�~X����3�m�$����ac�98VkS��������$��xTM6G�	$q��y�[���itČ,��wl�a8�f����H�`���Mn��Y�}���K��>����1�@�>�ң��������ąY	��k�Iפu���o!�̎�e]Y��H��D �������������4�s<)��樲���7' `��=����U�dO�͏H�o�����I�#P��-{#^}�M�v�t̡���ܱ(����d��R����y.�F9l�}�?%�/HG/�̯8�G�w�M�O���:�)=��X2�-�����A[HI�w���~�����F��ʎE�K\ߐ@�-�������8��	��z;�=K}��7T�:��j�yz��nb�n�H�{F���2h}J)E���/����4���{ܯ 鬒�Pj��z���ۥe���U�/�,R�,kH��X:{R�:l�JAۚ��8&��{�y�]�p5|�K��Pw��[�{u�1A��J
^�M3P�@)C�EI«W�q�����85�54�Rq 	y��n�J��*���-:�:S~�l6�������OQ�ْ�,lb��@�{��F-�\�	nͩo$�'D,xdKR.�J�
Ri��`tOh�&	�)@<
�X�uFeQ�sʆ#��(�/Ⱦ���\`$z�yI�U�l�^���A9�a|8���l:%��@&�/v�"C[p��,�[�����?-.�ӫe�:��n#�rO��0:��rH&,m��Q�����д>,�#S�6{�~Y<K���UX&��C~W=C����c����� �IBc�<u,kg��᫁�*�xX'+A_,M���A��ș��9IW�ȼ( ��m�.���(u!.�u��������i�>W*D���B¬u�0� g�ߠ��t
Eߨ��ҫ&L�=�������ë�q$���gN����2u�cCC P�l������♡��P���a��Һ�����j��)}v�ɍ�l�g��5K���T�I=GC��yL�|@�0g<?;+?�?�p�~�O��������هX�gT�)��	+��G�YP�ւ�aVX���2��`���'�}�=(��_�T]�a3M��w6/tkw#��`=v�7��ͨ�K����m�t'�ו8�>��ꮎ/����f��D2C�ΌM1���\�׆�S8D��P7!���'<����$ܸ�ק4�-7nu����S(�`��.Fd�����k�s��)�[��|ಈ�@��3���Iۖ�3,wP)�er��l��Sh���V��N�eKU$EӋ�;��ŀU��<���U�1x�w�Fgz��%�vmSQ���iY~��uIٌ�`���L�ٌ� SQB��2�����F�T���p�������2�~�W&eI�+^��inh)�:�E�AV�}h�63r�p�zf�q:�q�#'��6RCH�(0��#��Á	�d�oz��-�E�w�ȸ\�ȡZ5�c��w�dU��|�I�5v��\�v�� � �-D�E,=cC�i���6��'2Qq>L j&$K�:w3lٹ^��gO�u��KD��'��(5QKWē�*�?��}Si��@ϟ�Ŏ��O�d��2�b�$�w{O��8Z'ǥ<x1#��&Or��\�xă,��6F��38�^��J���C��ݒ5k��(^����Pi��� ˒.�h	9�~��k���M�5G�1�0���C>j�*A�a�WZީ�'�О����u�R;Se��5�~^;2��%�-{��e�.]�|8��`8��xr3�[?M� ^֘��uy�k�#-�T�a|ɗH�Y;$�3�(uvҏ�\���-K�~��͟�0\ ;9� ��*3��;��k�����pi�7�˟����N�F9��U����5���|�7��$s}_\s)�&�l�sm^;#{X༐�U�St��i��NMA}r�|��^s�r-햬���I��a�x^�GY��ђP{���=�����Y���^+�]Ϩ9YO�n8�رA6���1�l�p]�����D*J���9|4��D�h���9c��rW9��Y�ִ�L�������*.f�Y�-�X��X��_��{��ug�N�h�X�ȃ�׏�+�����R�s����2UQ��y2b��Xm�D��+�,sJ����!
�m��I�n8��s%,%E@�c����"�e�D`X@��
P<�X�����~�j(9�������n@� �ε�`�&U��*uߜ��G��=ү�#у����6+�f�}��?�{|���is�!2)IU��&�es�H�&6�˱o����fL6m���T�?#��dS���=V�@N�&>@8�`%��~2-w��w��#��|,Q��0�{�x�O��\#f���A��C��˭XdP�Vd.�V���=�
^��%�QQ�%��$�2������w�+�r��.ِ��e�j?�Rh8���`�{]��1�D�bbڜ�z���/2!�N�J�g�7��/��D�B�Ee�Gm�W�j��N�VNI��Z�!��� f
#v��\��Q����o6N@�Z�U��3wT�"� ��ND\>Q���k 6)-�/��j��Za'��tQA�H�_5��h'}�K d�亠��x
H�� ��]C��3�٪�XC�����'�c����|=�^�m���7�S�&�^o��(�d��_n�P���>>�,ș�4P>M��V���E��ν��k���M^�����T<�e�A�2w}�3��i��C�-,e����ԟ$��Z �cA~V0R]�^��LS��r
����V
�l��{tV��hS^`��u��'�	��0�<��<s`S�2w��륎7�"���8�i�Q�)$��m�f��E{�hc�]3�G3}��8
iy�����Ӻ�N�����|��)�.������S29���w���䑥��p� 9}b$���Ț�$�{�.|��=����]�����]�h�1K��cnџ۞��z�J�3�0tr��F�*h$� s��;=-�YRY䔧�8�����:D� a��SG<k�MfT��|�%�^C��!H�öv9M��s]��^G�� �ڛ��X�(��V��V�C�ǟɻ�����w��ZMe]��Xd ��h�a�!!�<6��S��6�;Nt��2J ���t�����D�)t���#K�8Ys&V-e��.��X=�E��u��\,O:�\!��t�s��CjW��u�h8J�D�-�K�dt'�"�QaR�w�Ϟ�aމ�:��]�M�N_��/��*#f%��g�A����O}��'�E�T3����a}8jQ��:vsS���E8�������L&��C�k-'��,J�p��1`�?��dk�m������%kh�Fq�6� �Wr1�+(A�!5�:��g?����ϖ��n%�/`�w�L���a�J���l�� `�&��)�:��&{f?Oj!�;:{�%4_=0�s��o�4) �+Ǣ4I�����W�CI.�L�M�*
���d�Y����j�w�ë@����A]ڍr���I���.��
�q\2�5ʤ.{�Wg��D������c����{����%�QM�'/8�^�~��T/�")�����>�zg[�OݣФ{�b�m��I�v�I�Y�.G�3=`.sث���V�l���IV�����~�!0��gQ��O�p�*���Y}��&�'��.q��&��y#�<|�y��.��i��(��{<8��w��<WF�-{�NP�����P�(�R%��ub��;�C�2�К�����cg����'X��7w�(��`4�l,�e� Bֺ��#��j�L������ӕ����qY����e����b��6�n ���#�kn���2lZK���,j2zQ"�u�ˮ+rT�)31M�_,ruSN0W���E�U���L�[EȷFɰɁ�y!�(��&��DD��Q�*l�k�WU�匢� 6�x�o��4��9����Dc.�&'���T�U���g��i�u����~�$�ȏy5���G�2Ϋ%�3C�m�!<߭/��z���f
��4��|�@�L=�M꬏&�v�X�%�c�^��$/�7{}��9YO�:aF������{�@x�s-��A��q����b��9��~��;�%�����N��Y�P�P�ڴ��e0x+�n�eЉ�h��;ǌe��ٺ�K�VO�ĺ�Љ�ޢ^Ōy�<�Z�������Q��˻�^$���N�6�J��s]
�$�e�^�Ђ����!\0�a ���m���[�����8�q�Rn��|��s�/0��͕`KS߃�$f.�8˹ۜpM)����P;7HUfHXcL�J3�8��1� fB�r�R:	�d޲��	'f�r�o,j/����R������gkC�f�V	A"�g�kC6_���Y�����	zr��s��e��떞VA�޲:���r�}j�/��w� A��a�L�MU*� +}�Q����ܯߺp
�S�}ep�5?b\�V���O��~�p�0$4��0]��zz�yo7s�b:Z�dRAV4�ìl�Yx����x�0f�5���'Ʊ���h�J�������<�'�u*��[g@
��O??�&A��k$h�[�~��j�9�W�p��'h���O�i(#^��-"�!�''~�TΝ�� �÷�����*�]I��TC�����s�������5��R*�ލ9�����Sߪ�n�
0Q^,���5����5My��tF5`ЍAnB�ex�%��Z�����#�$���E���b{�G��Wpf�n]��`��/G���ށ��Zaﺟk�g�g�e�����d�[f��fM�e�'Y���������5�s��)T�� p���V�v,��
@�I,�n�hv��e�q��������=>Ӓ ��K��Dt�镣�y,T9<4.̯X�Hb�)��E|��ǄlRee`=�	xӁ��]< ��l싯){d�rT�by��?$��W�΀��1�䝻]��n����3�����=�������� �S�����?�B��Wg��@f}���{�{"�}��rV	����w���PŹ/ok� X �f���s��B���#��	�R�8=�_b �uSRn�I��L�j��t���]Ճ+��3�G����v�ung`�Z� �
�C�gO��­�`�
�/��I�+��,�P���l��,S�~��	�Ɏj"w�0i_W�Ej��� �b�3߈�gq��l����Zb`� 5����4i�8�S�r?���X�ڀ���k��͍���=,�/j}3��J#hi}|����ޟ>��p��/^�&cdA`y���1�y�I^&�K��/��$`ʫ� \t3������{*bi�ؤ����$�##���0��z�lKBL|���u�5���'4�_^�\%G�2�];��sZ\�����m��A�G@�Z��C�0`_8����x��!��jF��p�yS����X��a}�@~y��۱�GJ��FaV��-�!�����,��LTd�+q������/`�r������a���E����TW%5j	Uf}��{�#*j�ֹ���1�L>y���W��ŭ8�������Wϭo&]�����.��������!���o����SO8���4�&V�,��iX�-Ř�`�J�#��~qg+��~8���gbU�akl�o��]��7��%J
r^r�����pɥ]a}Ϫ���Twi�����#b��	�}:u�u��Lv�� ����W6��<D}(2����#�����Ɨ���3���ck�B�!g���$U���{Ki�M2t��3��@Z��k�cC�_��	2���r�O�7�¤�DC4��N�6t'���p����H�����m��8�$���,�[V��2/�h�!�p���%�� �{�\/~'.�N�-��`fK�u	-��4��Z��ǆ<`Ev���BI!���$Ie���gT?����@���*fP��$�U8Ma�BL�z���� ��k�R�>�h�D�qgTi/<��/ �}�s
���{� ���é�Z��6�r=z����[�Q��Q��nF�W:y�l�^��mh���ɥ�4�4���^��M��S}&C�����:�8R|���3}�>6������jHyX�}tQH�7��	~g�����#;*Y,j֣
�R�g+�}e��D7�o&v�g�~�ֈEH@]�&�B���x��o������y�✅ATN�鰎5k������*,E6�3���
�åN�e��S�֖1�." J�������*Nɯ
A�G π�^=�T�+���چ�x<��&eQ�(�g�M�f�e����J��O�xTR-�3�U�>�9�h�+'-|뷂�!g��@���S"�0V�ΐ�O.�P�<t���I�=�3I8A��6?��Ց�U�^\�Wei4 j��Q�n6��Gӂ�n���4&;�}s�������� ^vy힁��l_2`�����K{+�51���`VU^�~��L�Y��j�$lg�>���  �q���k>�~�p��7h	)	��8��PZڂg^��}�M�� ��GE����œ�Y��9W����+H�G^�ٲ8S*+�Ԍ�䉓�rA�2c�(��E���}#ml���qK<io�g�$�V����{��pz���ȖoZ��=��Kh�OD�o�l�#�΢̆������m��C�X��&@����z��i&� �?�P�﨟�����k�Y5!���QK���\�`M��2�v�`�Վ�;���Гo��22ڧO7�{p�M�Q�<���nШ��/?W|y�C�[�5'�Å`��G�����v	$Y���B�e�WZ���`SC)�_�2�f`ůk&Q���X��rA��(D�Κ�=��A]XV�������+�U�\����`Ͷv��(F�1���;'�Ąm�[p�v��������%թ�I٠Vy��IV\?(L���n~��V�(sU�kױ1 �=1+nn�N?i�o�氄6�����i��jZ;����ۄ*�7譁�(x�M/��f]���w�AjVM�<� "�ZT׷1�p�	7�(�,C<v�;i�Ͷ5*��:��M�
�.�6��V�$�;���Ih�.��<����ޔ��F���}f��]E��l:��[��hY��07���+宺�J�۵A�y������v��R+h)�P�fov��&��N�J�oĒ|j�3)�<��ϫ��s*��Y�~�<����C��s]X����8��KO|�xzO*���C&��l��1?�w���vtdE�7�Ԟ��6᯺M S�"�ԖKO]Ȃ���Dl��+��S���ִX`V?��g3�p��;��ŀ�+��Fw�m<<���$db+g�?�(e2���lM�d�#�Q��MJ�*����[��� ~���f��Bi��e�̾�7�n�\�Ґ���i-�������46����Ɵ0@��f����v�|a�]�ǿ�� L��M�Z����ss^Y�L��~�oأ�^���;�]Ͳ�55[�b����	;�а�_/*o�N �!�ˁ�c*w��5]Y��Uw+������_��?hw.5|� f��������֪$J�N���I�a
q���rIᙯ�-t��P���,�ۣ*�7������/\��Θ*lC�{�0���5���@�xX1�g���@����,��w���v��qD���bt���<�N����|�#ʳ��C6�k<��~��_~Ag�j�'��(��V����4�X��xb�z��`�hU���Ϟhj`��a�q����y�A����7��@L�g�7�����^�R�X�R(�6��߸��gŗ5�U��L������d�7�}��"�Q��2����utw�R�x��ĳG�����MK���YM����XN�|�L�(�Z��lƮ]�z���K�*�~zpcY�Vp׀Q�c��t�ڤ.�~��]�ը�"1��;mIV��X�.�p�V.�(k�T��XiY����N����&1:ʰ!���Ir/��g@���y��j1��Ej��>���%�>��|6�.�l���:6W�}�+�o��
D�֑u�#em�<fM�0�?�K�y���'�,C��YhyI`����E��1��3�1��*dE3���´[z��� �$Fq���:|�u�=~�l���5}����,��k��P:W4�^���J��$g���
��>�"���)9�r��1l��?e����݋��늿O�f�� �,G�"v�i�ɥ!V��SϞr���	�.p^1�l������P��vԃ��=O�⢭h�*V��RN&O��r��:%�c�n#�d48j--�E�ŘG~r_�Q�H9��g�!d���{�. ���w.�0�#�!����r�+��� zՑ��,6z5E%��+fn�
���Wch�R��oSk��
jL�!s�I��-��`�a6APϥ�V�&$eLK&D�!:�jʈp@��*�}���ʱ����I1�%���X$Gr�d4��L�"�ٽ����|�g'}A�u�@�%Q?�u�-%^x�J�r���>���`�ɛ�[���[��Ez�ô2�13E=	���:*�ꚭ�%BY�0�0�E`�=�e��.*e�u2(��"к�,�2��̒�M��yv� ��<Xx�B�/��d�_���MiH%��y�״ȥ�*s�>�tM6�꫹�c@Q�A��&k���= a3Z0*ցD)�W\|
=m�Y�$��t�A!	S�6 B�E_�_�6��{Po�c ����.�g�N��¾��%��]�ů}�O;S-�ܶ���˨�Q�굵l�"���͹k3��V�(�c��?QFYf�R��x��`2�+V}�u�Ai��mBTC�rt�층�?O����\sTY����������̵b5�nyh�]#c���(��b*�+� �	�J���a���Q�����N�]�I���i3{�̰vݸ��H{��6�A�3ʰ��T�U�o�	�(ɝ����Y��]~��#�5"lG��X���L>���O�>'ӱWJ�$����d�@���X�����r2���}�m4~�ˀ��4���.IC������@:eN��F�N0��@��Ck|$�t���Z���e0;�`8!x��,P�݆ԛD��x{Uw�\�aP�'L6?ț�`��
z����)�q�!�`���&�x�A�~�e������;�ܠuע�/��G�*]�T�(X�B��%��]������Q5�[rϝ���5s����w�Tp�G���T�RZ拇�-��pѸ�#ڞeܺ��z�L��?y���c���6�eӀҦ��+��h�z-�d��*�8�2�&Kҙ���P���Э,��h�����Q�N`��]	v�Ԇ�Ey�{�Q���(��@~�`D)܄F��p.��`�� n��#W�fٱ�Q��_��->�;�`��ϖ�)���䟪�$Z�k�V\�������,��	8�������7�����pi���a�������MZ��$�6�.f���Y���,��lUx�����K��|A�3�P<$�<,�3������ۀ�b�T�ǻ��ϲB`m�,��&	0�Re��ݿ��/�,��;:�*\g�H��N�h|���@�ɸ5i��7h���rD�8΍�$��:��ږ��fa��0�1%�7�;��I�a��A���X�хi����/2)�WQ��g��E��]6vR�z+?�#�S2Hv����?�d�E_�,g�=�.^��RrEV�痠BX���V�zq9V���z;��q�O�f5N�0��5 �q�|]�� ���={y j��~0Ϗ��&�6}�^���+�Gy,w�<�7�4a7��VD��^�)��Y(r~[h��^S���[����X����p?Vg����6@Ϻy�ap���Q����{�,!=Z���1�����ׂቫ�1�OAb���]^~s�?$��G���'dS���c�pp�z�R�n��ڴq��ߚ�e�F�����(�6�����=nn�������>��22�be�D��ʳ�V+��V��_�tn����u���k1b^�:B)�#��x�V�7f�=�?	� cQ�Պ��E��=)z.'�%R�	!&��=�A��+}D �K4K�e���)�C��Gc?�:�:D��tԧC����1����8W�#'�Q��6Y^��Ο��7�*�:�5�LV��r� bỴ�B1p�6a*x�J[��k'|6�jML���H�X�d�e�r��؞�'bM�q滽]Sv)*#p%,fTr��~1͑چK�i���k���Ï�&g������E5�����lSS�7�Up�,����v%��g8�1���&h��cG\=��X�<�x��k��*��7��A��y>�3O*�=Y���<���
�~��k��)3_��T��Ή�f�}��#�kg7�vJ�bO�ܐ8�`j��w�;0?BS�D�h�H�0��6L�
+w�y�}ƫ݁B|��i�
(=���k�f5N�d;�/�`�x+���.��d�i��<�*�d"̒��m��˻_S�
1/֞us�_�7�lV�/�[Q5z��5���P�C�:���5X̝�Q@9)�&&n���7f��%���JI0̹�	-�m��9��E�9I'�y?8�z3�3��j���q�Qh�T 9�0���[J��\y3)���߃��C�t$��C8 �7�yJ����Ê��W��A����5�P1.��X�Rd�����S�Ϊl��xQ��0=�LΆ�otC����D��(P�������^��b��VP�-�/_��ڼ탽��3St��*W�th�.�hĵ�Z�D2�\|xtc�q~X� ����3k�p2,p&��&�y5�d�0��,�m�܇�z���_xyoԦY4-a�S)�|1Ш�l�X�,�C"V�2��
	`�$�%t3R�-{'��$&^�
��%P�#��qW!�U�5�8ӥZ��ݿq�]R�sf$`(�p��Sp�nڂ}�T�>:[�]�LӨeG��3�#�~�zgMx�)I����h��I�
��u��iWE�Ʒ>�Lo��5¸���_�c�צ�$�4����RM j�8����5Ҷ��9|��#�zr��W����p���J�����K�ڿ���� X��mR�6����s���]d��"��1 gT�WDC�,��10s#?qN��q�� �eI��2����u�U�'s~|\1�jly���,%���93JI�n<�x�#�_�qM�S��=GI^m]?|J�<�y��N���6���o�t�
�j���;\�b[����=���n�U�l�`kho봛�u~|=�?B��{�|��-��2��k�UB�7�6�O���Ey�򊓀c/8����f"���!J�� ϧn�&� #�,+Ԟ�1�9	P�j"SRi՛�8�O��ҿ'�C�T�H�q�U(�a^.���xT�g���{�����a,�I?&���T�u�;l�2����Pj]2���(����WsƎ�#��`>?3�����i-�[��h(�wc9ݘq��k��E@o�ٱ���E�i��bL>Z�?��{<-��!3ºDa�J��M��Y�-�K ���TO���%��lsRXcG~.v8'7����*
5��a������P�Q��T�}6�r��=�n2�?(q��z�����L��X���L7�?F,v)�ӷ���������'��1�b�K��z���e'�0��؍{�_,�!5�6����K�2���e�A�&��AWa���0���Q��I{}竷� ���v�����i���<�}~	��Ő�G�ܫĕ�F\ј���*M���^l,W=�a����c�]���)�����̺����Ypn�(ϛ�\Fp��*�Dҍ3�GH᷼޶���>���jϓ���)@sPn�5&�^'�Hs0>���h߶hV乃քk�p5R(�y��� �X\2,�]�ʣ~��v�"7�`���טͱ�ĉ��*٧���U7�TB�g�5h�&'�g\�4�9��ԳOSƅq���D�k P���p���&Ղ&�wKѻ$�ܒ�P)��)Ե���@gL�S��)EW J~\��N��V�0E'9�j�K_R^�\s���M(�i���$����3P��*���C���[��b8�G��j����=�2�@�/T�a)+IGI�����?\�g�f1U��mB�V�!q� �~�	��q��s��WZ�_��1T�ne���	�p�gb���[��z]4w�z29�ڼM��F��ud+|_8��F�\�Zt��NI�+n���(k_}f��O��j�3��o�)"�Y�0��z ?�9�&��?��!⻼�z�Ll��{=�l焠�����\b��g�RY�j"�� ��z��_�=���.}�<L\�Ж�Ss�,N�k���k�6>��b"���W;Nک6�}�oʸ�-#_D�@V����CY���Z\C�;#{Ohdg�T����CAȿ�s�l�.�<*x�� ��3�f�G������NQT��_֑/Ԣ��/W)��MBD��ڣ̮]�"�	�ƃB�����>�6�=����=� ���0�_�K�������hk�͂KU���!����=Ձ�e�ӓ+v�p&.:f{���M�sWcT|n���m�#�y˞�-/��"��_ā{m��s�EW�oD{���ݐA�h09�7?�U�� �ݰ��rϾJV�*�mAq��Ǿ� Jշ�)^:P� ��(J��m_�j�o�u��~e�*��Kf&��X�3%f�]Ҹ��^�q��}M�%P�K6�Y�mZ��-�2j�y9`��nX�}��{�����+�g�8�WÖ��E��~�k��J)�u=�(&o�t�(R�})����(	C^�7p����
df7�f$">���J=oI$�	�봾�N�YH�����2m�
��ho'�����֛YvE��Ǵ /=�����ҋm�Ld톜^��x���s��Z��
B���k���Mp����|$㘵�����S}{Q�
8 ^1^� �x񪳶f��-A	��<9��{ə����N�	pOV�LYL��`->&�������q��.pu�Zp71��w�8���wj�>j2u�(�!ЦI�\�G�!b��'���T�x_�g�8�1���D.*��/q�	�;����s�H$S�!U^""��AԴ~�j�P�͋�Ǘ۔q�Z�y����7˘#������(h�,�罋R���+��uLSD��ԫ^`jMN�
����ͣ�ˡ�le���9�jy�J���h��_~��ob��g_�Τ唘�RI2���FsA\���^J'ЇUZ6����Åu�T����oW7�>ೲ��m扭�L�hҨ���U	-��"��֫���;&�jk2����d�E,����b/)_f��q�S �h,�oMz�دs�8��lo���`�n�\%0q��vz�ϕSRIi@fpf�۞пAV��<�x��R��͜�-���o�=�[zD􏺥�f{o�n$o;�A�xx��C��cp��@�Jx��3[AtE��VX�l{��"$O77e�2���w[d���#4�>R�q����
,�57��)D��3|�x��aJ|h��ÏHi��iQ�#kb:�Hc�mʓ�mG9"���us�M$�,�Q13�ٖ�S���S�.8/q_�({h\�����Uq�}���[�	����&=�x�L�ȀF�N?�_0�J�[:"Z�t��$"�BL,�)̶e3S�R�C���}-�w=k$9^�>�́���I�����j���sU�t�:�YH����$�lmF�:ǎ]�u��C](���e��r�)�4={u����m�=�{Y撢[��y�q�N�=T�@��{Z�j%�c�&��K'[55�"f?��E#����N����%V�Z���M_�.�c�}�0K� ��/Ž�������AW=��8N�bhK7(��C����[V1��az.�Т��\��yqq�Mw�*�K!�!BC�\� 1�=^U�B��WN#}��ڟ������.v��r����q9CLjl\�q������h��9t�ɗ˴�X7'�h��p/TW���D���;}�UO�T7�<��qd�%Ky@����*��V(�A��s
]�O0.dG�HK�@�rFA߀�����tZlT�K���5>��Uf����ڂf��1�&�8�}���|��.�H��c�r�'xn�D,�jk�ƃ��FB��%�^����{�fG0^���R�}ǉ����S�A��t����y~sQz���iV;��Jh���&��*��~{��9�}�B@Ki��Asw�/h��|�:�	`�� {�����a�{���M�QK�����N����x^�(]��I�Q���"����W c��)����^o��>����a禥%��Ăt�Cŋ��~�������m9|v��*Z�<c8��E��9-�X�I���!��o�}u�:���TlT���,iv��נ�p��KYŘ�}�<;#�;�ϔi�܎b���DE��*l2u�gp���۫(>o'�4µI;@A<�g��5�c��^�^�
𮙙�;�������G�{ V���"N�&��g��;{l�F��0������&�|n��b	�@Q�o��Fcd�RL)[�P�%O�}�{�Be�~>��iz_`u=�j�s�T/�4Gw[����+�Sw;f��?�>	h4VpƓ�a;?���0A41X��t���-Ld��X=���J3'f��3�7����vv���	�!���B�0d!|��`eג�xΎ��O)�&�"-?�v�M|*��__�Z�.��B��43�n@��T'�JА�
l̎!�R3�8Xgϙ'ے��O����R�9�3a
����-
��,����Ӥ���9�	�+*�j�O�ai(�֭M0�\�d8��C��0赋)��<P�L�o^�DRxh��;b6D`?�:k��a���qZ)~G�����y҆y���sq#�-�*�/b�^��V؇J����ԜMb�k��i��9e�������,x�ۻ5���o�M[x��s&�����y"h�ad���4+�?+ D���?="���c?e��џ$֎>��p�<u��:Ǒi�2�wg��&Z�6Ʌ�}�-fͬ=L�j�w�k�al9-`1:�7~��<y-�Π�7��ї��5%l��P���|z2�,ߣi���Q b�8��}7���]���B�)�o��ϵ�ON��_,<GW����/������Iߪ��i�T,�e���3��Q�Y�`��]��7��8�h���3n.Uzr���Жs�I	�śP�i��gۿ�������Z$z��!���1�Ѱ���H�QO����(m9��`˶tx�f��2���=ƕq��D@��4|E!�+>���ً$ϯ�b�<{����rp�|������h�cU�׆p�MYr>��h����As�`�8쀲���8aJ�i�#��l?TC�Vf���u�,��bpvo$N,��ۨZ��u<��DL��ݦwX�^#'x�sՈ6�Dm��F�1�M�)�y[��b��]�?�L�7`�Q�=�93fBi=�#�-�ؼ��L}x��4T.m�x���ly�p����#iƳ1�m5�ỉ��� R�8�&R�Q�5c�1��QBh��-�m��]�����f���� �O�p��ш-|"-��b|y��+��������=��2X@Y��@�=�R.��c +����)GG��@dk���a�2���?��k�;��U9<�<M�n��d1��Z�c�7;�[�����=���b�陫RV�ys1�①�r�@e�^���^�(�Y���̈�m���^�H���I'eB\x�q�]MI�ǐ(zm�!�S����tv_�z�Ջ,,��>�W�l'Nͱ�\�����W��+(�%Jx�i�<j�h��"X��Af���4��GA}5f���iGC,KY'�Ub�u�S"g����[*m�Ի�xD�K^��y�c\�tE�j*!�Q"��[-�p����aW���{(�:�B��Tn� 0��&< ���Rg�I�|���X¶�X�
�'R�S0�e&Sk'�A<�w�M����g����3�%#t��'�]C*�G٨�~`Ʋ� E4���>e�q��S��=����0��.���JdĈTsz?�����F��������UW��ݏO��J��t���J�BP��o�7�����s��#EF��]�;Q��Hv�b���E�7�2�¹M���VxPT��r90զ�o�C�-ov��d����x����x��	8SȞ��;ה�]去�*fHZ�m'}�dǘ�Cm�$����+<)�k��7�Pu��HXr�� YΫ�iO���a�²�El�/���q�,�_���=�s�4��$������鳤��F~sko
�����#آI�L��5��PAC�"ꅧ�� �&a�6�{IuIl+y@',y��zs�|��5�P�G�!Ze��Cv��O��ޑȽ���^���QS�-R?]�f_|>/��h�&g���Ky�4�]yE�7�E����ӫ�\x�.��ݓ:��[�f 
�K?S	{w�.��-d@�
�R�"e߮�.Y�ҥ���iA�OJz�8?���#��5��J�p��#�1^�OMXe��x8�f!3/�UN��]��{Tn�Q����4��\������z���f%x��HZ
=A}���T�꬝�~�-U�k�W�����'G�^w�)s�a�W>3����ߩVta�ܴ���}���LR��5����k�q���x6�O��ן4�E����-�m�JD{&f��̂t�t��-�A.x݌|#�|쎙[���<��M@i[�0Ȱ�Z5�c&�'	���ʏ�]^��>��G+l�*�� 5��컮M�k�mʮ�/I��\Φ��� چ�i�P�A2��e�e
4��Xb�G�/{� &��$"�)O�@o��؄����e�T�:#jUd~���QTEA���iλ��
g���b��sb��ް���� �JV���S��d��\Lt��d���$�rj�\/���8�[Ƈ�::�$s�:N�pز��}	� �����F�z.����8G<@ڟ<�FF��,hN�P/O�,/9����+D���h��k?H�$5f<[0:O>��R�xڕ3��N�$�+��:H�Hp�D��_����8���*c0��&�˫�F��sdy�k0�+�c�oˆ����u�DjɊϼ��������ޚ�����
�z17_#�%��8/��ky�&ٓ�uMSF>bo9�s8`�q )f&�V��?}��q�=�j;�_�B�w�2�.tQ�`�չ�FŜֽmA��Tk!\�ڭ��f��%+ގ39��G�HV��� �#(,�Z����:r7&��U�x����Fo:7�,Gc��k�RJ�@����s%ϖH��y5
Q5%���i��'w��}��|�տ���]�C�b�e�ie���4<A���b�9�Q��Ż��xgwAA� ��nѩ�v0�!Wt����?s���<5��At�mf�J��1��7�U-�Tj�dV���;ؤ�|�6o��b�o�_Խ�b�D�w� yK]ۑ��*�r��]��CE?I��j��'8�39r�r)����������:���?M�>>�
z�ƭ;wL�}�O~�$4�w�6����9(r�v��G9#H�_*ɭRf�a�*:|��;�o_hV���=e��Bt쵯���P�${v�������#@&����#��'�E��������p�i�G�7�61��|ց�f�|�_=�;l��� �������\p�h4M�i!zG��**�I�n�"T��%�����ع�	��`��
&�38����%da�S�ٽ�e0P��Ϗ1�E�����K���+ߟ�� ���0З���N�ŹQW�a+��ڠ�Q?�e]Z� }��ÕE��W�L��T�Q93��g����U8�:�ߞ�^ԯ!@�]�(��KΑ�����v��S5޳+!8 #�j��0�<ӷ�s��9#�#ym�c�c��"Z���ոݓg�a��j������n6��/\��|�}Ʈ�VGޢ��0*����r	6�Ghߞ�����XRg�_�ly([����H&��)(��ڂ�RfQ�H�]6�)3�"��i�=孵#7��(��@Y����	��_��E�F��B��̳A �h?�e/:R��R��M��7$׎��J����Mw�֒O7��
n#d(��h~�ק��%���A��K	 ���N݄Y�5��Q��N3��7�I��N�h����?�K��h�B�q����q�S��v�G;C���.����ghϓ���g��Sϯ�Qh�1rW@᯷G}��oζ�c"6��a΢��&�%枿��>��D�:���J�GS�s�T�::�5��ėC'"j@�S �2�٢�[����$4)2�Zy���6��eb)'�1X�N��rO�.7��̢#Q�[�Q9�(�i_�T!'3�j�T� �EFЧ��3\��zƶ���T�0�[0SţX���<�����-aAR|ΘO;���I����������f�'N?3Au�:*Rc.}��kv���\~��j���\i�!3ϖx碕F�=���?�Mn���`��ƀ�w�ǋVJ��+`�]��UR~h���s�eD(JE&^$��(�L��N2C&�v�p���jC���%�؃vY
'>�Oi���X��4�C�N�NQ=�(�!�q������\n]�havY���!r�ϓ��=�p���2�v��yuS1obJ�����1Nvu^��G/�ԯ�H�;�jKY:[2X����_+���g.���`�U��V���+<�8ȩ�+��MW���G_޶%�`o�=C��xj�&� �R�����h.zn�Gz�i�8�$�Q�k�G�����'?���%~:v)fSZa��h�}w��%��Wb ހMX��{sA�+�V��V<iמ����Y�b[~����%�1�W�r��RsQ�F�찷�ZH�����+���"���1(�No�0�����g4ҽW���N8�ё�x�y��ܴ+	¶-����{RdJ+�� �#
��|����YlX4d��Br1�Q(qd^e9 �������t�)#B��[���y�,r6��[�b��u����;�-�k|4� 
xU�E��,�a��$�t.i
�? ����;q��r_�`/ѳ|>�D�u�"Q�D�#��%��d�\M�����#�th ��g|���8���ʍ�%1nK[�)h05QCP!x�0��"��@�l�H�.ȍ��zn?mK�� c�P�8�J9��z��oP�8��g�,b�N��F:�.,��:cde�� N��Ao;�)�9�7�}�ʱ�
~�������v b�I��?fg�, t}�N'o�HDi(�^IV����(����1�y�y'����Lx��b���"�B�tm��^2��H���xZG��q!�|�%޹�eb��bS���[x
-�E�lY�4�K!���5"" J�5���;&��2�[Y���n���H��{�6Ʋ�NC�wEݬ��C_t�k��9CNP��z�m�*�d@���ޓO�&��;�;�q?�����l�t{I(�ZA����x��&1�B%�k��f��GKX;#�m]6J������p5��\������t�f�J�c��P#���!I�XOb�SHZn��P<u�c�Ӟ�T+�n:n�U���t�L�wf,��|��M^QЈ7�����k��Wr�0���F \�nc����l�D:7�g�E#��,.� wfn������kґq��'s�r�
y|b��
���]��O.A�Mh���3� 9t�A�f�W6���s�jC�<�4{Vt��h�]2�SFQpmjv�O�Q3�@������/�}���~à-|�՚�z
�t|dʧk��ވ�W���%DĬ�AB���	�+�j��n��?��������)�g��<<vmP��B�0�`��Z�)�s�[5�W)�����-pĠUdC�ßk��p�e�B�ҵ��B�_�A�b�8΄s8���Pc�Df�|�/��X�C������ђ-�A��2y�	%�]ܡ�A�9O��Bˁv�\Ы�ݹ��W��"�-N��s9j��
S ����iX�Z�"��e�C;BZ%0\U��&d���!0�Si���(A	
��̈́w�I;$�Z��������`:����`���������_(Q�N]q�:��M�"�-{��zL�O��ýrB�/x�����(˷�E�����cQ._�.��¯Ȕ~�yT���`��Z���r2S�$@M+]�n�F�O�P�䟩���@��,]~�W��<J�Ǵ��lhN���q��ׁ�<KC�6�e��D�`LII����׽^�6M���.��޾$hR�鍹Yq�DEڒ�PGJ�?�}|�L�~�yΰ�ݜg��tn���1��iO�������)��"�^��H��9�l������:��VH���n;�&�a���K�?v������TG��6ѯ�F�@m�P��R�2P�R�t&�)~4J���@Mp��15'T,��`@3n
ÒG�|���^2}*���"P����*lcl�}F(z�X��5C$��JK��>��ZLc�W�k��}��V�JZ�L.�{���{�w�,�?�4�5l�(�5e6/<�U���=�{V;ta���i�O��W���Ja��ͪ�b��MzO�Q��^+g�4Y�:I`boM�r�$�H��h�x�g�cR��r�������I�U������ѩK(\���s��>A��\�@�q?� `�d�$jP��NL`��ɴ��)�4郺���L�RX�'�ٔ/6�Z��E����!���չr�x ��M�g��H��y�����rc�h@}K��ހ��}(�Ċ�7m�� A��2-�5I�|�x�솵����nfbv�}����鳎u��B;�t�wB��h\5�H�2��-�	א����ZGzì՟�j;�#B�Lě�>�D� � �e^�m�t�8]�cyE���5�|�.��� N^"�g$�y��sm���k���*ǝ��u��R��%��[
��ʎǧ��l|`F��H�I��>�H��[�o*��i/�P.�Z��Ӄ/ښ�z�"��5Lq�H���K#{� ����2�  ��t��K:�ME�B}B�e�]�}q������m��rB�^h$��++..)�zn��q|ۈs���ͥ��S�AZ�v69����,���S��Z�,>���a8����0n����P�>��o }2��x�1�w#��Կ{���k	-����������Kh�z�,��m��֌�a�,�tnb�w� �.@$Y�UaX��r\x5�1+�fն�ާ�A�ۿ�W�%�Js�$k�1����Z#�!�8��E~���h��T
Z=6<l�a�q �U�}��DQ�7$�I�`gi���(�t��b��s���U4�#%۰[5�zq߇�iX��pr$	l��N��z���$ޛ�@3�0���f@���OC�Ɉ]��l �Ѹ�22K�n���t��ݙ�������b;�5_p�R#���yBow�����ڿ3�b�����;��^�>��dW��C�u6�pg��y/_�2�ן����Źfp^W�cB:g�#2��5w���Vyc�8ׯ�82ۺi��1B��_�E^�ם�G�<`">z�䁚�PˊE��ʤ4�A�K�����s�����k4������UɃz��O�b6{�?m& �/U��Z�~�[C.^�f�v���:�AM`H?װ�'�����lep�C�G��k��G9��͉6����h��(>�-�ϩ�V,�k�f�ŮS�I!i�t��,&I�f��f���O'V��D骐>uy��Dj��)�%��g�^7��1?�ϕ������uL��l;o/@ό���@�*��n��%u�FC�� ������dȫ]݀�zH���
wz�-z��M2�Ҋ-Z5����4�0���n--M{��ླp�f*�aar���H���ll]Lv��.����F�䳮���=e%�wc[̗�-�f>��?��{y��>H�>6T���(�g%�����%#��a�ht�C�35~���Uq��$�y��Sv$� ��R��S��Y�L[ŕC�(Bi�����6�4���`�O1,	t�RW�!�R��	�������#���f��+�Q �;��|�͆uh�������S���|�8E��`-TC�&�tN�3J������+}\�yP�Tz��>�[ǹ�#���[��}H�J���Az��d-h�=��R(AJ��\-*�(V�`&�Y�ѐl_�g��#��ݺOO絈$�lV��:����3��πL�Ю�fHK ��!�&
w5�a��nB;Mи'��j�?Ȣ�Μ�C�QA��t؇#w8W
���]CKʬR*�`V�{��_�ek��#��I��HD������ft�3��[�j�0K[X��TfO`�h6U�+��7P�ށD�A|���29�k���꭯M�]X����L�Ŝ���Pɘ�UXM������*�1]\}ITȝ��2ǽEC�O�D����+��̪��e�t9G]�/�MT�s��������`ޞ�l�D�1�@��m[�W���IM� I�
�=�.�L�.��7�/�'�v�E�l�9�&�ljl1���F3�W�ʗz٠W��N��p�(ŝ=|@}����K��s���ֻ�.lo��C4 ���x�k��A;m%�}#�ׅ�bU`���̒����kZ;�W�F�6��
��/��X�y���ٳɚ���U�.pl���&KO�EK��Aq��c�k)D��p���:�Ҁ��'*B�9��I���7ؓ���e���0K핿N����a 1���3�_��oD��>����O��*�e�fk��H*+<��Y?���|���e�8��'��W�����m���.�HYE���F�ռ ��j�,ɫ�_z��O_�X4��������
H�]���ض��7U��3Z�˽��޸{{&?b�μ*���7��q8g60q-KHu�؇�C�q˚�:��0~LP�H�ݠP��DOÍ}��A=Caku�ި,��s-���żCԠai�`,rw.`��I��>�q��2��s�<�����]:�1�J����x-�]��N `�b.f�B�޼�?����QS�\r�~O����-�w�t�"2~��P�Nv�
� �>���ES`��>%�r ���K��w���^~
�]����q�����h,0tܶ�)62U�E����MG(���E�k�!�P�%����y�?ϳ���ڃ���ܧ��D�q���j����*�Dͩ�����S��/��K=����D��0B�4��)bf��Q�@*��b��Uu�s05�k��{h����V֠= ��Ɇ*k��ˆ�,h;���.���*?��_�Μ�GIap��H ������>�b�8Ȫ!��gK���ׯ�����5SeO���I[�P��8�N���7HF�f:�i��R&Z��5����*-���weWPX�l����[Nz|��[�"�.��%�˥'�t��c�����si���D�;�B-WƜ�E݋$jicư��ntR���6�l�V\�/�W-2��ߜ �Z�n�|%���H:OD��!ъ'!/Z���k`�G���\.�u��~�l7W\k�L���Xt��>�#�\�JFض\�w��D�$1����?��}�U 0Ac�5���"˰�S��Cf}qF1[Z��|��M�K��eP�\�$��qs�R��PRC���r���-���5����(�A�u���E�Ȓ���j{��� ��z���u�X���F�c|.9�_�j�A`]�����Ӫ����i�/Q�}Y����AwD��	����<�6�4#���o�v[�:���?�h,2=���`��@�O����b��^*�f�(�~}��Fu;X�uȥ_+��ƿ�)�ϫO�����i���X����,nOuY}�6[�~]\�MA��dGd�$�%E��Q68��y.��2�Q
��x�
;~�fc�b=�:<�X	�=��?����ů�'��IIKs�>�w�8��&�m�X���v)��	�������V'��
�5@����.'�F�j۹���H���MԞ�����L��Я�(Oa~M�e�c�E��ZJ�"�&X?�OC�ti�˿�X�]���]h��`;���H.�[�ܶqX�7��LVr�W�ag��+��C0Ψ<7/q�:�ٹz/��p�W�Q]1�\��S�_$?����V��O�<���8�_�~
k�6��4�8���BS2I*�L4�y�@��ۻ\'v���
pN��ŝ4ӵ�k=3��%���&p�����H�6��k�!lk����u}��Чb��r&�R��i�B���m�Fw*'>Ɋ�IQ��j(C+`D\T�`���:���h�W���6�e^�*��?T�<m�W�R5��8����%$�N+��˖�B ��)h��T�#����1��<�ȏ�b��}���8&� bỪ�[�#��-�?����/Q*��=�ᔕ�f�P��j ��޾��-��[�^
��#s4���	�6�!��1���`���>܉�����v!���_��@�B\#���>�S*U�M��ʗ�&ۿ�r1��3�N����6�D��y��쀚�S�3�fb<�F�O�O8i �4P&�������I��4>s�~ό����C��p�/�=�g����3��:����f��[~R+
��
�a=�O	�5m�A�?�p-5��M��'eS#.g3w6��6@�����⛰����)$מ�r�[�-� �]f]���O����ّ�J����)n���6�v#"���*|��6�n�n��bzK~j3�F�y|���m.{ Ȭ2k3R��I��f�u�is�rY��.(C���ɳ��ەT���?&<�j	�8$�I����c��#BZs�6�4�c�A�'�^?�3/2<����E�+U�:�2�x�V�w���A��+�o1c�ۅg��W_B�JlQ[s1\���!#q!��$�('���N+1Q�P%1�4�kG�i��p�/��̗a������r�AQ9H.1�J`���"F��~���,����p5�ܸ�S���?,�d#��ތ��(*.�2�	H��/�
�F�Y C�Q���Y��kaOA�3�w�a��) ������rB+���NJ��g��p�H$?~J��g|+��V*��tĹ����
�P�jvĻ<�ZV��WC���PhI4��Lۥ6��5޵���7�'3�-젮Y2ӏ�{�ƻ:�?͔��#��G��	��KE8�� Q���7џ���-�����"0���\#T&Q;�)��Z3���k��,o*�mi
#��7n���PG�2yW3ʩXDg�u�⺃��W�(�M[+��u�<o��ވ7�"a 'p�nu�zx~=]ٜ{��+嗀�w��b���Gg�EH����ɵij�Euw�̘M�0����������ce��t�[-C���6���n�o�D�^�^���_g�H>��f&�Vk��+����c���6#��9��)"e˜���T*�-P�F�zV�;�ki�gH����8�����8zh~R��H��gd�]!�����X?U����=�x�`�Q�xU^`$'�����?�P���=O& �,ƚ�ĸ᠃f[=��ec(�����'�D�WP��-��6�*��>��؝�F��e!�[��
��%�:�
�z��`Y�wiH� ��;�}8�R6L�a㺲���Ʌ�%�t.&�;b��E��b`�|b��Q��nI�i牮�k|b�n�|�"3�_O�j�(�3���x�jj���ǰ���.�á;:Z7�O���Y�I#�9!%+�kb��V�!�o03��=��1O��/��\�q#�N��N�&��QbL��1�c�%�f�TbR�_�)��������6�L�כ|�SO/أ�o���Մ]�HCz{5Oq��%�{r Q����ц�ܝ�M�dyEʞ5��9!FM�:��pJ�p>|�*�A�j�t��W����a+_V��]�'9m��� ��셰�1�-XJM� �T�IQ���B�p����z�33Æ�i�����Y��Ɩ�	�#��%��P�G��_?��S���?#��!.�RS�?_
����ԣ�j~��U+�S�3�o����3sRnD�Ͳ�9�&���#�>��}
$�e���I�Kz�����5B��$ r��U�&��7�Sщu�*-�ӅE|�`�����iL�㈆�.!��O3K��l�'&0fCژ��� �d�pÙI�����@��4�ƍ����yl7�֠Eӄ�沮��9�SyòՓIҫ["o�(����Ay�f��xT��p��V�c�0�[�/Tl�ܠ����e���Ń�r��NXW�)�
)g8���&�3M�	\�	��j�c��w��7�P�ë+�Ã|9K���8+��a,�ڮ*�Z4q;nX�ǟ4�Č82A/[)�36+���np�&�q���Q����K�@���`�zJ�p��~��ϙ�%E�J��4����D����K46��\#ǯ���mԀ	E�O���G����6i�m9�a�Q
��$�},m�\�TT4��i�YW] ���D��n��b����SeiACY�)mE�6�ǈ|����&̃�U���]ܖ���F����6yu�Z9�q:}��Or~&��/�-�<�@2̍� ˕��y�U�����T;�+�C+�x_�Nj����\�4�k�5n����G�]}����FC��~�f�)�V��M��v��e�mV�	���M����a.����Jl�C,���p�~��c覵��:�i����7��Ӂ�k@�d�1G�y*:fN���V����?�:���_Ē�~�H�n��g�]���s��v)������M8�c�����r�Z਒�^���6g�+�p�?�9�h�DƐ�溥w� �>Mmܮ��[������2e�JF��׉��3�����N�9	�BSr�J�2b�٥	𖭢�
�-��8�>�� Gê�z=<�9���w��M��@"d�Ν�:�F�Ҽ�a܂�*Z�K��5�bZN?佻o���rǗU��E���k�M)�1 ��#>O�3�l��.�Z�#&���k_WӋߧ��j�̤�1���,�r2����Fл���J5�.���S#�B�{�XR�;�>�+fT�*I�K�'0ܒ#��P�i�Wi�ǱA��u�,� ��v<u3��E(�F#��ˎ/�?��٠&��c��*��,W�:Ꮫ��b�j�̉�$�T)��*Q��.p\�&aPεr���p�4*�e�z���A��<K�p�GʤF�'��&3�;ý�\F�}�����A�K��p7�KW�-�+��������37�x(S���ҍ��C4�����V�PN�Ӟt�� 5RH�d*:�GU�F�>Vex�B#j��g�w�t�8��i79<L����"ƤZ+"H��b���cK�W��a�uarG������ϥ>L&�u��	�1��E�Գ,��ׇ�޹?����<AmQk�y�&�`:�yw�]��Ujc�{� �ɜ�B9nW��������	`@sV8s;1� 'FOv���}N�w�t�x���Du6S���y��k�d@��X�yDe��X�t�#��w��8/��^�7\�U��f��� �ve?�NW�m,=MZ�o����F�WwqT�+���*� ]��=�������\��!�6����WE�r�0Br��pz�aԢm�(=F��r��jX�� �=������}�r�3<�U����`�K�K������!��bDD�ץϫ�o�?�Gv����H�1�����0�P���`�s1��YI
��1���0Y��00��a�ՔTdg�r=f�f�<|h��'�f�-�V�E�c�:U���1ޡ��܁�|�Ea��RJ|X�Xb�>�RD��U&c�}a-Cri��כg��g�^"\f���Kb��_-]�{���J=v)0��Qjͦ>��6�
�����Qt�@�Z�`W�n�G뾑�,����k�]��$z������9�;�oW��4A)2ga�������w70�W*hc1@%��_�j� �Mmu�w`��h��ϔ�O�#{;ꈗ<�'��޸ڸ���нA�b,4H��ΰpb���'���)�Օ돔���.7��,�Ϯ�))�LG��k�W3-W��h0N���2���J��e�@�n��k�k��?�����aҕ���ή��D�+�2dSHAJ�Lb�YC�Q����'��N'O��=l�T�_u�L'_hX`nJ�/,��˦��c��\��G���M������ʠ,^o�w@����Tu���k˥�dg8�q dwxxY�*�����F��@Yc����Μ}�V�)��?���I�Y���=7Ö�?�4��h˧�6���^�/>q�z���o�\�8A�/G,��O9��aP��QӘ`Ў���%�	�� Q|�5)��-O�+�w%Wo6�E4p������9~���Szm��.̆���r�p��]�>���C���F��?J
�&tM⁔���
�E��S9Xur�G�tR"Q�8n`�����P��81�Vlu�ؑ��'k�&nL�L�� ����1�^L5@��� �[$Zf����&����*ҍ��.މ��F�8���� ��.�˨�"b(���\��w���ę��0��K��(+�TN+�	�.�啽��ރ�p>q��~���PF{<�C�FB^�L$c���_�y�$��1�Fܟ\1����%̄1�r�\�>�A=pP��0{��g��UX� ��c43s���6�������%�/����#a%_���"@W�L�f�z�a�`�5���zm4|��S���}g�x�-tU��>cX�(s�z;���e���O���u!dPX����Y_�t(ˍ���E�
�A�M,W䡌��a=��u���Bk>�
����=U��o�A�����1KN��%ز2���/���ĺy�2���i�/'#X�j�Y� ]�nZ�m4$��=�5�z���8�oD���,^��*y
�{��(�2/�Cv���xF�-i�rgJ��.\
�7�_8&���>p���k�\�DC#�����sW	�;��v(����34ﰚ��tl����Ai�N0�8��˂�l��ϵ���_�"X����	(u�0!f���v��
�/`�"��"<�i�U3�}(�q���BL0�Z��|)?qpˀ�Uw�!��'���\���,1A��5�����p@O���_�((�VC��<���#Z�D�`�B�����v����2�~��$��#��0���S@~/��ē�;�n�!��v�%(�M��R�6�cN����1�\7��C-�%�R��7I	�C
5a�S��vMw�&��EJ����XO��`5� t�5�g���1�5KE4?�G�]�􊅩�U���]�i'8�-QJe!���z6�9�Ud���^X�1����[d��f��5���ƶ3b�<H��N�-=�r�cx���(	���σ��m�@~�MDXO��U��.����V���t夸'6�9�������PC���ha�`|���XiįG����6TOx���s��J�E*h�@̎�{'�@�}�����ug����mEp�K�#��kzY)|"M��*<�N�0�Q��J�~q����o(+����8*?������`�An�+&�9��V��e�Ԩo�f���r��h~��s�]���q�e�ߍȞ��F`�s�j�-z��(@���aE�/������^�P�_����b�F�NR
Wv�T/����l˼� ��\6h�w�ry���#�]�%Ҧ!R�He�ќa]ꈠ�,�B���Ց�Xt ryv�h�Co>|ε�d���O���J����ivxXH�wЄ��=�Y�}�0�fH(���b���_	E�?��Cùo�ӑ�����tڤ-d������gcqV��"�c��ۺ�{��n�s��Yq&K�K��:��0ۣ���ejx�9Lj�@B<�>I�a������o�@��+�ó$���s-�F�n1Z��̊g�=(:J�lyL�79�k]P�����VIASO�>=�񣑇� ��_v�TQ��A���2�֪���T���
�0�3�q���P�5�!���+BA��EV�2��P���]$lg�u׹Ťт&�x��L��U�`>S��B�-��0��$���r��x���ذO���$����}�\%�gq8݈�b:n�KqŞin.�G�1�;�K*��}&���D!�H�3����{�\�|��a��p.���7��62n���m1qR8��l9�I�h�M/Y�S����@���)��acZ�,N) �ʡ�`ho�l�D歵<��P?e�̆{��x�)|@�us���d��z�WƑ���E?\���13o�����8<�����V*	\яHTc����Np�8}�k˜eHGa$���jW@�5W�YC��5׌>�;�%r�z�o�����Hf��َ9&�n)s���L䴃�f�T�%�R��?��z9L﫡,a,�7��zZm���������Mhp[�\����z6�Z��B��g��Ht7��A�י�Wd�Pb�d� ���Δ�j����SwKV��He���_� ˝N(�~9���Y�V��I}����pw��`�>k򤂥jh���*��?��l���ZO�.�uP�z�K��R��e�ߥH�ݫnԮ���װ�ýo42���*͒y5B��_s��l����[u�D�B�m�����w��V�p�F�wɂ5��F�^���ܡr�QC)73�3<��^���֬��HƢ�+���1���Ci8���,)r|!���<T�L��$���AqD�T5Gƹ�z̦*�W��N%z:ݵ�i�n\h��f�-�I�� ��bY����3�����'2�YvL����$5a�G�+L�_؈U?�6����:�P_C�䔶&�^��M�Jl'�6i��4�P]�˳���>���z�#�u(�)#��U岗~���u��Ĥ��D��Y����fp�`�u�R1�NOw�"�ؔ�9�eP�u�(g���XS`0��໱.J?��f�����Tz��lh50�h 4Y�h������@���S�]��s�a�J�YW==?ؙ�b������Y>�^����Y��S���128�w�"�7Dw�	JT-T��r�eЍx�w�8�wBl��j3|�����9v~|�;V�~��y�k�0b9F�Aѓ��w���K�� �+�36t��)�:�e���*�<E�]͊���Ŷ\�e��՟����kC��̒�3��������{8�	�Mת�� �! �|V����)��c�P Sw�g�z�u���Z��G�tSs��P�JA9z�ԫw��Lo�?��� 
S�E�ti�l�6��u.�~zl0sJή�^h�)�i����\C	�Q?%k}u��,{�]�"2�e,v�������)$�N,p(�8�\�)�|���YȯQ�`��y՟l������ Z_7��ׂ��g)����_ː���judP��0��_e�s��^RA���"׍�p�z��ԞދG#�'}����3S�(�翲���U�j�м�؁�&�~ *xdƗT�_��B�m#)�و�e{'��*�������i[
���3q's������UA���Á�u}�A������,�8�3�-?��K���Ξ�M�b�p6!��-s@�p�SX|mS�x�c��>��Z�A*�n�n
����YNxVL*��h��~��s�T5՝�ˋ���6��W�	��!@9'���e1\_��o��¬M��k<Yo�{O*�
�^V��SN%_:N�����qw�T�I��ӓd���9�5%�J՘���,:����u��]h�;��NF�e�X}xmN��f��M	�)��L�Lv�u�p$�V��a8ć�JX��n�b�1!)1���Vpљ*��8*�F�}o��3�[�^��oZ���E&�1�0s�rB���bäSdr;6Ǵy��bY};[c�Sz��0p���A�i��f�iVm�~[�Y��02B�֕��j�*�[d�f)y
PB���C�5Y�	�]`�[���Z:�^����{48�>�t$ע8\��*>:�:�����8�j��<��R�Ԏ��m	|�Fn�aΙ���p�0�Q�8�C](��0���J[>�������/+ U�='yz,������>T�p`^퐓!�ڨ������ҥW���R�@/;�f�k��B^l�1V�e��h/���
���$�d$fY	
;��.�I������r�i;Y�ͫ��k���g�$���9���>��V6E��BOܸ����!�S���0�G�)�B������~�04"�L���$4�i�<e���l<�G�'���Rd;��!��V����ֹ���#�C�vF��~{��*q��:wU��,��dtxe���G�r�M͢��o�iQ��p�tV��.�;�@�x���M]�6��S��u�B5#�맸��mOQ��dV�Wnɡq�3�w�u�#f"YF�8��׼YǇ�Kw{g�����$������ut㛣iuc��>�pˬ���!TS;7�M����^�و���,��'���VxKɪ9<�<"z]�Jm-T�ʏ�uu�	�#��b �<�0�xЁ��������	�x�[VL�*A0�կ�zl���˅�7?���u��X
���*�?��)��|6�<��X��(%ç������d
=�s������#�*|T������G%��VAt=�&$^�#�D|N�7��	��,#xhx���y*������x+v�C�@��K�U�`�ug�����*uL1��O,~}|W$�F�h?<�Im¯(n�^F�(7;���Od��±;��#[�; ٿ�%�Q���cBf��p���$�ֹDѮ����H�N�����7��e%z�&
�*MQ�vA���Aِ��l�.���#�3�o좪1%Gۊ���k6����>x�-�(1*v>8�檣�nڠ$�T&����j�� 9S9�w�s�
*u��*�B�ңM����e�?I��k{�,��8��x�ˊp]<8ɔ-W�n�zK}qG~��w�R��'�Ya�N��e�:�A��9�֐��;��� ����[_+��v7x	������a�d6��������o��������w-5v���oz�Z+Sլ�d���Ln	%{D��J�< �1tе=Fi��B?���{�^�C��F����+��i��V��F��8����}��fL��N�����p{"u��T��?eQ����~R|ލmt^��ۜ�LL�9�&rkCD�rx��p�����!�E�z$j��q����I�(�uQ}�
!>/�f-8:g' _W�j�j*����fd����}�~���l6���x�`e!��l�[.ս*���D���q_�)H�����7g��Uz�Nt?����	H�%���̎�ND���֘V+S�\��Hg����>����2�^�������g���1�i��S�x.=G<�0�ωL�(�l�qB��׋ف�펔N�(|���1�6?z�%������H�2�	]�R.0��Ma��Z�c�@0'PW�9�en�vOUС��C�u��J�a\�{�'�2�{����>*��ї��I8���A7.�|��/R����ll�|q/��,�p_�T�%rL���XZ�i92;8��^��brh6�[�J !��	�]B>��[���lz�NI�� Ϯ(C�D�����h�TP�<wN$e֐����)_�ɝ�_���l�4ic]�S�S?�K�6z����e�3�"'��dԞ'�*=	�g���N~�Z���fgX�m��p��#i��	31��$����-R����l���`�&$=bj�R�ƫp�ِ'���t�u�e:Qǜ���3{���Z�`���-޾͕�pg��1`ѻ������|�?����tԂ7����a	5JD�,�i�P���i���d{�fK�	|��|�D�����iK�������EȒY���q�"���~$\ӑ��/� �{ v������+`8է�wGza�p;��	i���_�bkN�,��xm=�R�+J�\,�:�Tg�f���K�ˈ��[<�}'�W�D�7�jV��%�޿�-����b3�~F0j��OԕUXF���1mn�����ߪ������[�͹�,b���^�:�U��9wor�����8���'g`u��s����zX������N�H�(lR�[.�ݴѩ:�Y�Ŏ�y��V��|�g� ��ܑ�^�±��U=?kܬ��
��)˺7m��jo�����{�F(��̌�T9'��w� �Z"D����t�oW��èXB�&5^W�{�N�:3\2��=PLxױ��7���	����� ��-D+�*ښ���P��{��[����)�ܪ� �#ԥ�[�`~�j�J �̩�}�f�	�M������{����z�T�b�|q�������̲�T���2clM��B<oߟ�'�rhfWxoN=�Y>�G⻯����ev��-�x0��!2�p�!��X�T����[f��Ae��!KP��^TtT؃��	����Ú�#��7Ig<�Y��-�	�a��� �$r ���*m�8����}������^`>�#K�+��#1�� tq�ݐ6vbh�0b�,i���6�����[[N��[y�O_&�����`][�0(ƥ����9��8B+�����&v�v�Z��UHg��d�ut�΄����ҳ>G -���Z��G������h�������(�h1��4
=�P���x��>��4<Z{���L�}�+%� ���xj2<�#t ��5Dm�yc�G�4�T�pX�G��Mm�U�y�:��kW_!8kqQ<S߿�m��i���!N-�\��o��<m<Ks��m�)����D #A^y��'�J������I9�����m6��9R�$��0.�`; �I�����m�Av�� ҲZkǣ�c"�@����z���얯[H��U'b�AjΓ��'�_��F���ۆ
X=���b@��yX�udV�B��f+_�xg����+�^
�2��6�VS����"qb~���]�RبvƘ�����t��#Ʌ~�ʩnb�mv�[!|��kN�7���������#	���"��1p��JW��Q�|\��i��y��5���t]B��F�)��d����ǈ��Su�q��kg~eW5O����-�d�/�	�1���9'��݃�+�g=�Y�e	���a��B�k4 �Aj�$����~��9c�O�m����R��ه��<j�њ����zͽO�z�^5�0�ݹ*�@T&p2�V��;U#WL�usU�#�Кc�$�;
��m����'v��T�����&#�,{����i���X��oa�٤#�,�+��	����?R��+��m���l�Py��!ڣ(ӏn_m.K�9��֢ ]����d�V�$��Y�(��L]%� Y��]e�-��M�͖�+�C�g�I�*߳m�Mk�6!=�������ށ����*yTV�"�.g1e�m�IzKm���^�EBh
�H� |Ҩ�N<��݉)T�4E8�z>w� ���&�7�c��<�q5f	�p�����_���9��Y�ˁ%����H�؎��|�v���g��o�5б�����?ľ&�TU�� d�Vh��[��>� �
��!��P�]n�gpFx�.�C!�x�[.(MΣ$Ō����A������)(W��F��ٮ�8��Ϳ݊��l^r�O��r-�O&@�c`��Xr��\��VM��]W�?�8w[��n���y��W�?xX`\4-N��:��-=��ǀ=�x���O��Y�� �}R*���zޕV:u� ��_%<��:nzx5_�t�#����/����cwO�-J����\SM�uC
�`�-xvc#������<��et�7�s�PT՗���`�g��7]����*�iAͮ���'Z������0�-�{�Q$�zL�P���A;on�k����
D���G��y���y���q�[W��]����g>q{:��]M��4#�1��3PJO�ىI-҆����o==b�u@�mSN�|2�� `Fu�#�ĳp�@�b�W�zU�㍶�w�<X 'iQ$��|�2���9 >ܻS�s'�.|6���|����$�	��`���9!'�I�5BnXA9�<��c��-�b���������Y�����_!�jb	���hN���FqH�N���vlBگ��Aq�m�/����Tw���B=� �	��b~/���n����!/r�CY���-��c;6����X���A�;��?=�i6'�p����r�v�4'K��	e�<Ko�=�R0�(f�6 �����֘���dsq�k�(5�E � ��V�;T���1~;"��E�A�W�a��m��L_�i�ɱ�(�*|����^�΋��)�A���?�w�5�@f�
�%_��@(Ԓf��Ď��%�|�:7Cر�k����UXM�Ƈ��ˆ�bWfC,1��b\������&s��0���x��Pĥ&�~�F��qCzX~��V���m�����nb�n댑��㆏�e���� �:ӑ��G6�;��8��/��J<�h,��M�/�E�R.m]v��]a���x��026;�O��o���a��8��B�[2Q̳8K�hc)�8W�l��9:����
7�6�#��i����V��[�p�� ����_�a��,ܱ���� T�Sc2K�)�647y����tft\o�}��`l{��)�u�m���Gv�a{���I�#���0�Z��U��J{�~j�ٶ��m��6�U(h��r�	�=&�_�|_%)�Z�����%�G�����gO�Ƭ��z�FD&٭X�Ѱ9|T�2�b�[ȳ�rbț/��NאG��,_=�/\=n�����Erlk��>X���	��O������G��H���a5��ԍw����]�њvj�*���@E_��/�L��y��*�Q�.�).4�PW�e��\V\�Q�v>�\�~���j^��"߱|��s�τ+�t���CÿHޜ��s9^�[�� e��h���u�bNqߥ��
���oAX{j�c���M�*��ثG����gK�wq�]N1�l	��E������݆�M��}�v��&��ץ�H��.��n-�:�tª�j��[;��pÛ�Мewj6�	Qᓨ����򇔤]��x��;.����۩��fZ!��ǭ�#���d��8�'�ɫ�h/T1�w3�I�5Dy	��~���v�L$�S	Iʵ�kJ���u�/$ꇾ�EEi�ʆ1ٕ/C�kT v�bKuh[���g��ph�V�
�˄��#�J��'��?|�X{L8�HO��\���c��7�SB��ۣڼA_~J�-����x�7�B�y�����``�Cv)�Ec�� ��,L�\�[y�0��;�P�d�ll�G�{׸}-L������(���zQY@�i�����(|��cp����eWg�!�(C|�A>����u3\��Y��Pd!�W?$�%�J��Y���ng$kv�<�\��?���p!�G��nR�������d��`�8;�.��u"����%[o�BJۭu�a<�qV#��`	��\�G^�?-�h!H���j�^���<�Ϥ�T��b�W�7�ޭ@�1�Vc�m��I�S�k�_3���2���} �����ǵ8B��B�X60��l@؆�)8�G�	�r�!Y��x�K�Zdڟ9ۄ����</����Ў?,���ݥ�1&]�ә�KH��|y
gպ��7�?NyQP�T��������ܕƏ�0y��+�fQ�z!�mءq��c�s,/{Im���3Wv�dq�w|��f$���D|����v�!��~�c?ѳ�
��ȯM��1?h;�y*��w�e'�F$|W�5��V�=�H�c�~R�x����@&�߆�'{{38ԟ�����;��҄�+�/sl,��I_����G�B`S>j`�����UĥYuɥ�5%x���1`z~��/�%�&��F/3����qq�ɾ�4ޜ\]9���:� "��?jޯf���.���D��?�ڃ��Ģ�������PL��Ϋ%瘈hA����v���N��S�ƨ��f�C
����H���C��ǥ�,n`�&l[�?��N-8rEPz��y�mFh��?|������t(?/?��`�yM��ޮ\�y;)�ˠG�ٻ�����LL>�)�	R�:�4���� j�����cߜ�]6O�����cZ���.i��(��S�Hi�P�ה��_����5�a�����A���:�V�Ѝ�%�/l��3�֡�{{6S�UN4��z��4�L �6UA�/*�o������n��R������hw����Zd��A�`�7��~�1G����#��\Pv�p��.~���vL���b�F���Jh�)B[����\��zʯO��j��W�5/C��|�h��v�"@�OJ<��Î��%��&̛���)�m��и�0����W,��*op��S���[�ݣ(6,�����'�`�/gR{s:�JC���������鯖��%D���ҭ��h���qlz1�4��u8�H�Z���i�Jf}A�)��K���U���ϱ��b+�IVZ���r-�'"��#�@���A!�TT�
��8�d+0F��gB�'����E�.������"){Ɯ�D�&���Pg��u��g9<�!cN�N�	�m��%�aSpϒʫ8�u�[T���K�p����aU[�,�'#�9��\'���T��5��`�(#�x�:&��#f�!S��5�ƴ�J��AF8oS�����J�g����GTbv�Mm=ERd� *�bG�DO�T��{�Y��a`b��l�¿��O�ħ��C
�ʋ��nq
��R�VYL�!}����-}l,�M����ia*������^2��k5{5.�y�,�p�hhZ^rC���A�!��;��0��?��#�BD���d�� ����(.��P�4����"2���,.��M�B^�V|��.Th؛TR����b:`x}��p�UU>~��T��� ~�/m�-�N�`��Z��&�m�9�j�%Ȭ�&��كi��krW���-�,�j����v��ze�?���nS �6�r:�ղ��,ۅ�'�S%����qn�yT�B�8w:ߺ�FSz�8��P�H��6�ө��8�z$�=g#J܊�yeV����Z��Q�'�����9b�f(l)������Aңj���VQ�B��0��[~܇���y�=Y��P�Z/�'�x،����l��������`�s`��@8nﭗ���SIp��.�;�=���D>P�9�)��ߡޝs[u��pp��'��LYC���<\1�U�Qࠐ�%c�,��]2m�U�xE��B6�(F*PE�Dܴ���F&��c�~ɹW.�9o3
6���\8JZ^4ԋ�iL�� c_@`.n��\���Á�У5p����Tf��p���p+<�^!�/u3\��bu��oKU �����6��o�^���|�gU ��)EoSς�W<�҃�pҾ�"�[H�&,L��Rk%F�9g���%�Z������=�X�V�/���3���Ց�+�&U/[�`��2�Д���쑯X��@��H�R��I9�U�1P�	���l^[�[�0e����q���Q��߫e�S��P7��@�wĵ�j��..,$�A_*�L�	����k�*�+�.l����I68�*nH0m�ɰiw/�@-,
�����w��i��ш�߉;C,c]@ՁO�W��"�J}�}���2|��"�WyHg�+z�����-,�$$�P�Э.?6�ҵm�@5�e�3������Ռo��;W�):sF$еw��sF��u���^��[�o�4V�<�A�Ʉ�A��$�$�`1o#4"��uקW�1FZ���"җ���|c�(�Au���A��� E)%�	�:�9����ߕ�#��H�yz�Ҭ=����I+���r����rs_���D�*�1H�)<�N�u�0��zv����5�p�³������[�7aLd'5μ�f�U�(Ԯl��W�τ!	�ǹ�#�2��46�,�bt����( � �p���-����CI)�7��4զ��	��u6mZW#� d�0���4*�m�\L��5V .J鶇7��8��O�6a)�B-7E��r��Կ��}!���;]ϻZi�0Kӆ����9���*���y����X��r�Oj��|�;Ml&PjkH���35Wߟq<m�&;�ހ\�_ƞ�� ���3:���nrVf���R�re�5��I6:ګ.�v�N���~m��ɪ�EݱuU��FA(`��U�'��T1/ڄz�d��5��[C����%�����	�u���Ӌ7���ڼ�o(��n�x�$��/��E��k�����E��4/�E�t׳��o<*=�ɴ�$�i۠� Q�?m�����8�^�:�g m:����.��c�kjPn*Vz�(�<���d�����׌�ӧ����ͭ14�;@U�O���d�A�-��T���&C�S͖�B�/]�v�!�5	�)��NU�P�����r�x�ґ�rG���$G�h�Z�X��0��_Կ+�3�I���R�y��ve�!�#	�%HMx;��S����c5�<{���U�}���y�����>�۳����0��)R~�hܘ.�Z��)Ia\���$����/jLjy�>p#W���bd��c�l���+�#� '�U$��eT�cwR�DՊ]��<T�[
��y��٬��C��w@�J��A�־�~~4Ps���!��]�:Ş�H���N�V����-*5YE�t��
Fx�����,Z���L���SߊJbD^yV-��fr���"W�DGi��:�_����6�����c��k==��9Hy�^Ո�V⌟ ԰hW�s�-�ڪhR@��|�bd����S`�M�-�v�쁐�0�	4���}�1�4��@ź�i��s���`�����K��c��	���O`0��l�Ĩ-p��.(�'�^����<M������,%���0-Id̮"mDH�^cvxD� ��ؠ��(�sw�e^jK�S�('gg0��]�m7���~�������N�sX�)���S��d�{(Ew�j>��^��*����_@���m��m�=$kʴn�%�һ�R�_%K�v)v�ds��"X�����޳f���c��UF�>/�𭌟��|Nq��L�Vf������l}C(V���m��/.<�0+�(�E�'}���hE���C���q��@<2Ք|��6ټ1���'�o}j�8pQu>�/x��!���)]*��˻�veҐ��6����$��mL�ܧ�����$ڶ�
��0�� �
��aW�mz��rw�~��S�;�'���gB�k>Ǖ|�T֠qj`�x�7�eo�~����}�o�m��cO#G����~��"{y_T8����*�s����Y3�D�����8;,W`��]�X�ȼz`�369[)9ׂ��@\��H4"2��K�ZZk���|�|ѝ���6>x�BP<��t��5KN�� �/�;x���⨬Q�X1ME�b����ϴ� o������rI�!\`4�������E����-�(Wƌ��m�ڤ$+�$���P�l�jOrc9�,3Y��"���'0)@�S�� >t@®��Xv�F�ɔ��Ȗs#[WQv�P��	��h+��β�kZW���۱��_�U�L^�$z	�{�T��yh
%H@w����Ĺq��O��c�4�#G�X��׳�<�:0	drX����̵����)�ͅh�a���_�'S6����=	��Ў��+�l�#�u�p�3���)Db2��:�R�>��K/�b�+f�@T���(��uBR���(��	�}�=+�Hx2���շ\�엟L�\6SJm`lL����K��X��P��^'g�*%*A���d(�Q3�A�3|Y�_��室q�U�}r�DJ?r7�;�=\{�gh>Q]k���A�#��¤���N`�C	�H���*]��ۡ�h��}I�26ߏ��r��������gZN233�L������ΕJ���T�d�z�������]�n��3�o�q���Bl��M]`C���:�zD�)x*ZU�w�8�`C%uש:Il���*���NU<>1�c�8^	+p���pC#hf�@eS"e�/^�y��a^�����եu�d���pݖg���Z�`�]�ڠ����ڡU�)�m���h�(�`�����m2���Q�H\8efڵ�:v=ѣq!�J��j<��|�A@��E���z��`sfO��W�r"��-}vLa��+�}j;7!}x�g�������Bi|՞�c�c;	H*gBLp"a�*�ce�#�mXg��ެ��n���D!l�ü���W����J��M��9-o3�rJ� �(`R��%�3��#VE��l�����/�ei$��Ⱥ�rlk��r�kn������T��dXmyT�uqn]��'چu��Y�]�3����c���w��
�Aߗ����b]��#��ݦ\���^�z!ܬ"�b�-���ј}T0�O����R�SGa0ě����#&�D��$�v�JRC�h�i$����L��%�QD�%ed�5ڱ�Zޒ[x��`�c�/�ҷh>�°�Ұ�4��� �Pi�[����0$#
��UC`+��Ŋ�n��!�E:��U�\K����p.��?���lt}���=e��7i���~�)-&�K��@��!����H�t���]�^fd�%� ���	�{��v�|)T���*c�-�gOi�ً6�14۹S�Ǧ>�V��߇�. ��3*c�k��i�β3���!���5S� �@O#Y���/좼���kHEL�ν��!�v�F��;z��2y^�.P�ڌM�4��c�Õ�(���������FHc�;%>ފ֪��V����]ta�&c��=�U-�Hi��ٷ��.�<g��A�h��£�LM`��5�l�\�gy ����n�K��>ڊ��rj؊v�H{rz�N$f{��,�,�T�V�������&4��e�w���ZYWS��|mlj�Vg_V��Epf���B���cKK
a0�����TǕ����*���drHcPf<��>o�r������U�*��(Q�$8�@d!�
�pJ��x�	3��V�-����-?P���}g��x���,æ*��)4��i����.��A�ܥ�Sa��8l�F��&-Vq�.8�]8{��@!f�^FO�C��{IX�6g�ٹ��.-'o�LC2T������m�h��4�U�ٌ��䠭*�Aw�%��9I5y'���
�9`�˖���p�5[��>�V��z����s�̒�9��[���#����UC:����C����s� ����+a����"���� ���p!b�m �4#j@�W��(z(�I���AS�m-ߎ�O`��I�ղ>Dp�
���v3�����м���E�^ù3p���fi��*6���������U7���8Q�su�wܖ���Y�l�1�/ +7�␲�p�Ns��A�(y��f|E�Ĩ���|�ۋs;Ƥɼ�t(p���{@����
g��$�Z6==��}/��
�?� ��Q�In���J�BG�]C�y��u`
��rLMf$ �������a��1lQ7��oh�2�_aS�a�4�ۆ�����)b�[vd�e��b��1:�֐^2U��`��u���b��P��k	U B�����)���7��(¼.bSH��B�Ռ#��R�C ���!�m�/�wA�#݃�su�&:����=s�5��d�H.�:�h�'绞}J?%���v�� iR}�d�?��-�8�o$,�������6i���֘b��J�T�.��w����&�ڧ>"Jӌ� N�����ɓ���ؾ͸�~:���C>�)�!�B����$��?�C"�%nwШ����㚻O�\��6v+; z�!da�+0�$��Q���.��H��?T�o5����C�O,^_8y$��;T�jSr۽+5��Fml�,������ J��5c���J����=�}m|�0���Y�Q+Ǉ�8Y�JZ�.�����K�v�@	
��6FUHj���Ɍa��w�3���Q��j�hQ� �N�����7�fF�'��N��s��b�T�"�Z�Sι@1�A���4J%7T�ԫz"�l�D�;�%��>XJ}�����.�g��$�ֆ��I�C�'���J8��N����{�dX��&��=LֵIY�H̄���_$����q_��	�l�`���!���!��L5�y���5�7�g�6�Ef3{�i��9� !��.������QtZ�K��T����M�=�gj���k�|����Z5���,����V�o�?�$���!2�ٺ�]f&Y(6��F�U�`��:G��:�I�;T�s�reuKF2�.C��s\�[Qb���������Fb⬶�P�~�OXLC��
����I���eS3+C����=�(}`U<��>
gR<9�K5~�y�>
<��gU�g��8�˨�H3��,c���i}�E�X}YMl����;��sm����}��T.g���SxY-��eDD�,fY�@���L�Bp}bS���_��ɻB��I}A���_	'�ԉ��  ���30JH�.�S*g�N!P�04h�۳D>�ŸƗZ��R�*�e��
{����BA+_ڤ���U���8��2�d���U�īD�K�Q�Ȅ��#������f�F���~ܝq�Ÿ-wD������ݬ��NU*�96��;��Dނ4�L���8)�= �(�S�b�w�e�U��Q�bB�Y*��Q��[�����ߩ9�i�6n�}%���M�13���E�Ԙ���Wq�Ơ?� �*U�bffZ �w��%fo�#�����P��UHH������J�E�x5}U�ٴ�}�����A��;Ob�)b�~������U޿HX�9')�n��9G���P?����w���G�$�oA-��a�a(X3��7��a�F��g�e��"�;��F%�C>���i��GP�C�y���\?HΤ���rֲ���jTvR9Y��Ae��4P�0���]�d`R�AY<��7=�98K��8� }�����^�y�~����A6J��7����}����s ����]j�cO�[+���#��{�
����K���	���ce&f#л���9,<:��L�ϝtG#���77�D֜ux�xٛ���	}<����N��'zU��g�Ǣ���=
��q� <#�����m�	][c�sOǑ�ook{�;a�����I\�A4<���8������ zս�[�c�����C.>��2�2����D��]-�Dcs]��8{ ��iT��1�RW�&�~�i��dd�"tk��6�y���a���=�Z���b�;7V��c_��;�яyԴDE�Ct�&�M�T����5�EN?�F�Rq�X��ӱ������V�F�tr�N�(��h�p�z���E�M:a���T�w%�Ů�U���*�d��ɢە$B��I=s֐E�ă��� Q7��+$Nr�r7;_<�a������j�/�R9w!;�R!Y*�S�Te�z��'g ����;}*-�ʂ2
 q|v�.-3	N�j3<�:��[�D����2@1'�? ��-3욑<^�"�����$����۔��?;\�5����}�B�Vέ�XY ��ian�5�݃{�A��\pJ٥-����i�|%f8ݜ�t����elE)y7ۉ���$�,�~(�zN��qR���[��V��&� ť�k�
��+�bK��&�.)DY�0ķ̙ ?��^�4�/�fP/�h�yo��i���0��a�}�b��F-2��RC�� ,B�cq���d��X���_JA�xsa��"��m��(^!�k,�1�k[����6�hɗ6�p��(F;�4*ՠ%�KY�O5��8ڲӲT9�{w��j��������"YAb!;ؗk�=~2ӄ��2�/8���,��_P}���G�I�=9���˰1;�m�j�י�G���%I� =��}5�s�L^�%�M��ۉD����w1+~E.�q�]�����?�����^�{7���;��r�rJ� Z��*k�Йq�}R�3keOe����0��D���Q@�v� q� ���.we�󚎢���3�T�>l?.~GQ��c�!aFp���	���2�ܪ�=����J���8�Y[Z�\5$�E$[�]����I� 9h�63��ˑ���G7��L=��F-�M�b�Ї�Ub���t��
1��0�ӕ[�KZ�Q_�K��F{�U��s��	�]'��ܪ�`�f4�[��=�[*�";e�p$Yu��τ���Q]������^�F	��X�D�IQ�zǨ�u��N���V��ӛ�/KW����|i8����1���*9�*U�SpF�{mISj��X���_����BѸx�7�Cu��~da�Ƥ[9/�\3!�W"L�C/�w�#���um8#x������
�LS��*��ك�(0恂�����Մb�WbD`��f���u���G ��~�}@K酲���uVw���"b����y/�G�a�'d���8Y�F��Me�=ŏ����vQ[<��Q|��k��E3e�uٖR@9q}9�K Z8���	Й�w�-��r�Q�}��u�V����'�_n�"!�'� �|�2g4Բcy�˲����b76D~�B$Lak���($»�[�S��dO�)��īs k�9�2�N���\�4��Qe����j(�;�gt+}%���]�pAһYd�A�l���=�[���-s��TJ��'�^LIX
}���DE;SvbA��O��ܰ�xL��K�I��v	��;1E�"�bM�$��}ڡ򐤹���>��+P1XA���W��}rҗ��p�u�1|fG����"o�
Th<3�����1������0�7Ϳ��"����S��U ��[|���R�1���V\�ʾXL!~a�
�f��i��!A��oL��_��I����A��*�Z���D4xTC-ʼ�XC���z� ��[]:K£�D-J���ϕ獽>�.du��fR۬� ��6N֒�?9����fC��rwu��>�ǤZr��}�<�ĵyJ��+�W���C�y��(ȼ��9w8��f49ϖ�n4v4l;��+xt�VM���
ȫ�f\�P@92�O/p�1'����Vyjr�� '�����$�&\a&ȈUI60#�@���N$����rr�w���5$J�X�j\k��$���n��W�����yx��iz�z�u���݄'!��IW�P%���y�������j�o7�\`߀ɦN\�n�,�K�&m{X����G_�Q"F�{Bv�(O��E��k�$C���j���l'D���f9�/:T�6�t�-8mɤ�!9�wV�;G_m�y����uTX�x��L�DkR��Ҫ O����������K��H��$zY�a�!���g�a���{�s���k��Q&�%=It@�6)���r�NdC��1`1Y�0�Hr$1�O�N�X]���K2uZI�� �K�eZ|��L�����,���(�O�ӟ(�p�N7c���!�4���2�U�8In^c�h�$4y)	a18H���n;�EA����f={'��]��6�����q@h�0cϤs�Oi�>�Ύku�Ջ|*�X�66��P��S�U��ҽ�b�Լ�y�T�Z|R���ni\<�U.]�Om@J�n������-6h��1G1�c8�&�h��7�A)�u��71L?G�}��!��M�47P�~y����f`}�3�h�V��&�����a�ܑ�1L�Fƭ�p]H0�=�{F8O)�r�EVs[,)m*w-<���@/�^�-3�m�Q����cض����C�W�4S���MW!n�Hk��ƿ�UIJl�N��l<�eMR]F��W��(
�R��*ڭl�EPN���~{�E�Y���+@��Y�T{�Pl~b�˸ۗ��=(Z=\�m���.N=��	w�;z�[�̧��"����yC�ى'Z����xj}&�pZMw�_���Q)ji�5���Y/�k٨C�}'�A���9j�̑�E�k���M0h��Ë��Dߦ��TƕJ{n
'b�?}w�P�(dȉ�v��8w[n��pK��'$���"o%v��_�5�p��ϸD�Y�u~��O��e�W��_1��`����ެ�.er���B�l0]b�4g�(��e�gT��ِ�(�wma�.6"I?iR��{	3J�D�G51�N��b5��?`䈔	)�xT$�b\�V�'s|Tww�!��&��y&*�D����"j��?�߂H��ož�NVyAs�ugRj��h�Xk�;� `�Gi�/7��7��k+8:p���g�$
��cε(�_� 	w�1(K��OpƔ=���	��OŸTs��Q\��~=B{(xB�������}����E�I�UA��^�n�! �<Q� �Cf$iDk�����A��`yD��K����7�t��»���}-c�E�������?�w0M�H�_��n;��X��ƚ����R���+��=����+�E��.�b?x	�iA{F?,m�|;7$;a)q��:�M@��{���"��[�x[洯�j�]\��kS_������gZ	ſ��8*xV�۬���2.3V@�)��p�Q{|��pOQ@؟�� ���G.�BSIB�msB7�չ���u�;�M� L~*x��=�&jr���*o��V���M���	=�3�je���0<���P%Ү�>�g����t�5�x|��P� ���Svg �ƓB>2'�L�CN��K�ܔ��\n�Z��^���l���ӺV{VfT��x��qY֎���"lc<�s�)σu*����oJV�X����5�����3mG�L5^Q��?W�-����֛���zJ�G�duR��!��R(�Y�D�1`<�˺Y̶��Fw�0ݭB��,m@����ok;W���O���Ġ��������nt=t�ymόl�+�b�TZ1��(�#f+W�cq��	���x�a.i������3dg̔�6\c�5z%NpKd鞭2��5���
4�۩K�R�4��wPï��xL�����1��,������A\Yo�i��%��hs [��s��W����>@!��M7*�_�x1��@�EiN�����~��>�I��`6�
�,҈8��0E}�F�P^t��u��X��J�k�3�P�˟%��M�_2@�����L�=���Y5vO�x�zT)�?`��`C�	�a�
����3�b�K�YK����a��X<�%��#�n�W2�I��FAz�A�0���>���h�0U,H;��Ȭe���/{���Y�U<�(�j�hW$ȇ�iܴ��V,��"n�ӃL|k��]��\�co[����9D���ge���*����T$�)�d��^�o�zg/*x	�-�׽ކ ���gB0h��'���I
���`	�o���X��f�ѝ�J䁤eb��J&<��h�1���	�I�*+�� �3U1�y?�@�@Ʀ��9��vӫ���?/�_�^H�Ƈw���&)!a1R�{�i���4��	�gpf��A��R�҂����nh>U��A=��aU�%Q����Q���_��2�I�1BQ��� �\�O��%]�y-*��Ef���B:�؎����ڍ��L&�U�;�"�(���RH��;�%"*L~��6���F 0�,� T�,��eV<{������Љ��H��%��}[���)y�O*�P��L��aE��c?t���P����z�(���?]giu��;̌�A20Y�,U���l��g���
��F�`��
mJ��Xvy���afRF��=���-w���*0
��x�<�U�z�ٹT�]��Ǖak��Y��
�I|�J������ȵ\�$�5B���>����Dw���v�Y)���%F��&K4�:Pv�����R�S�6���Bm�=rDT���\��^I4ne�t ��]@P���U��0�n�_�s����v��ْjyN���a
�kX����% S2��YbzΑ���+�g�A��<���u�om��`U�NI,Ou�	� ���QR�!����c?~o�I8��0P%�N7�f�^LMۡN6�AS�f�k`�9��1<<8,����U(���	�����Osb��Ӂ0=�{񳼃�9N�D�C)�C.uE'�ب�.N�f��D�Y�Ȟ�i
�8
?�`Ykؓ��%�����q�I?�5�~���^�`ORCQ��(�����<�$�� R�Sw��$,�`�ħsɅd�}��x����yu-x�"��N!Ct��9����`+z�pC; ��5 �S��uL�y�GDqǭ��s�-s�"1A�DDF(r[5ϯ��ˠ��;��͗��D8���p��	Q�\���*\�}�R|el���RW�&m�Ԛ�2.��p�[%gu����f�7pr�dR?#|��׿������ "ϴ;:�*ne�	�a4��%|퉆���m�N`�!Q \{m�Х� ��z���N�[�l�r�[;��s�	D�T�L�7��W�lu9�#j����]�S�a�k��FCa���z(�T���E��|�l��wy��c���u��n���Y���2���e2��E�F��n�Oi1�'����-X���>JX�O#DOV'5�:\�D��A��M	����C�!U�����E���>5%#�o>����)\zY��Os��L/}k����%�%�iLY ��0�^�	�=g�%fG���=`
DʂQ�l���o�r���^�{�����1./3�o��n]1>��TQ���0����g���E�4� ut"i{z�N���������w+����.�}d��l"n]�`���kY]B��K�M��p6��dx c&���7�q��	h��!{��~����4n��n��� s�����3e�!�P-�稾~�k*��`��i�YCzV,���n;['�M�i^����X�;�2n�\ ��溰<�}�j_�e��
6 �딽H}���JZ`��Yr�Os#�bǣ:�ڐ�Gf��b�%Z�ƿ�b"{H0�a���L���}��S^X�Y0g��0ު*0�23w(ka/򙻒=Z���3 ���d*j�+"y�~592M4�:����Q%����t�ct	�F��tD.�l��a�+�ޥco	*���OX!������ˠ�[��v�%+t�.��Z΃�Sh�x�$׺���i=��_N� �=4��.�Y�
ѱQ�o돲8�HQ[tm�pP(^Mۚ��{^�梈���C��}RM��v2��9�+:+5�@��<z7�TT�jGhLV��EOL���g)��)l}MQ����M%7�9׾�M����s"Ѡ=qo&qU�5�1�(�\ <�b����Oe$���*�I瞳�=�PA�C�0
"�Ӧ>�R��r!��3�-��9�o�ѕѸQ(��6+�m��j��÷�P�'��2M-}+��Y�� ��m����a�s'�F�m`օ�P�E���s�^��l�.��K�е�������H�RH���ގ�o#׭���,�Gw�>�KF�r'ςuE�Uh�$f�d̫���Y��w��n�/��ЇW�㒄���Tb����d��\�{�E�ƢD�G��'�h>����\܉��Q~��yi�=�����n#�#ܣɢ�Y���2^Hr�"<��(��%P���e�avl��i��fXQ7�	;�	M��z�Ņ��s[�_�v��q��cpV�m���[�O"4Z\YD�3u�[I���Ƙ�&����:���  8��sf�6�(^��<f��m�%Y�����ꖣULčo�MDs����go�+��	}��O��6;ڧ�9T_�h��^@�$kD�Қg����]�����/�
��O�S�pȉ��Iv�g_�M������z�i�:ko�wls�a��3�����c��B�	)�wXx{������ء!k=o�4 r!��Q4� �}܆CҢXv|=E�ގY�[35s=��t��U���ha�zK�\���7쎿�W�:�?d����O"J�0"mi��O,�^'SA�!�S�n(�#��ݲzf����e�~u�#$B�Hq��x'0���h�O�yR07u�#���V��"!�O��	z���[e�R��Fց���f`EqZ��u�Uc�\�~�)	q�)��u䶓�E pb��"x��J���h�~�z0�\/�PY�S~1:]�{/O�X�h	���N x��V��#%�׾qu���C!E���S
AM������C*�����Q�����M�	=�����9<c��I�ZS�x�]j���en�������G�G�)�́�i�h���,wG*j����D���)%xش�O��X~�cUR���%H��T�꽕'���}J��K�auG�m}_?�Ћ̭���dTf�ݦ��� a�ų�0�#^4t�F�u{?�F�	�5�ݤ`d�����KmȚ��iiG�+��}?�xS�����Y�B��f<����Q��w_i&���x��*�+ÿY�:,�q�U[�
��R6O!��t�fiK�k,]���虨���}1u�ǔ�}��"���1����ls�7wZd���OȝԯmZF7s	R�xt�2f D2��|6P�[�I=�]55���zz���o��kظ_Q�rߙ�6(Q8�:�6� �����E�&��Lޘ��E�W]��ٗ�'�@�;���*ރB��_�B��=9��R���z�]���^ϼg��b68���x�	���" t72�\*}��^�2��kN�}���}l��oc��ȁ�0U��|)�k�1E�my��9�'����J�B����_�+2P�2���è_��*���İ�	@����@�9K:�a��"����.>ެ��͡>8�j�=��m5��j�S�(A�<N���{/��\��FL#�ݟ���ث����#	A�z{��'�QAb���}����< ����B������k^�c��gB֝��K��[|\�;LBS|(������7*���9�,`A��$(�e�3v	��������c��s�d2s�̠�V����BfAwL`�? �Yf�W��	��l���T(���C�3qlD��0*5d��Ћ�7���!���X�>�In#PK��ȉ]4�x/]�O��
�Yx��yJca� �\	��g�u��\ķ��a����k# �3Tn�g�Fę��p�N�io�ŭ�������G�z��-!���IO���{"�ʣ��'�zل���<�}��WʛLo7Nl)��E���M�,`Kt��~f ַE@���x���(7L�N��w���ʥ*G��.$��OD1A��C1�����;,��9�D8t��#�T%� �@޴Ń��k�'���@��8G�;Lk�O�����ڽ(Q�-�XY[n�(��ȓ�Mq�ST������v3��R?��++�n�*͵a@�9��ހ8b�� i�B9˛��d��0DW���MH�(1\�/(�0`v��%��������A�rR԰ܜ�@����$	��bL�jku�ƻ+��ݡ�!@�T*�*�ǸB}��\��'otI~S}s+`(`�:�TT�_Dp:��-�X+�_����H�ts����}�z�GX}���y�H�G?k�OŖl@�״ȕ@���zH�LA�dH	��	j��s�4����v��c3���J���:$�	�f殾^ܡ�;����~K����]G�VbY���`s��,2��4jr�	��~��i H�VJW�2�?�kw��>4�Ǎ�����G���
�+�sGH�9E�ĹCo�w��$皺Y^�Y�W�D�{��#>TN8�L���@�~�%�k�ўt�C\�%�wc`}�������׽WK
���_��{�Ң#�9@�d3�m��j��|:8
b������\ ��-l=��CQG1_D�?��$�4��t4��)��׼�I��,��u�>�U�C��8 �]p�[R�5��+�;����c�og\�S�ͧ�%}��ˀ�ҷ�E�;�.t�|�f���1���a� =�d͑��Ȁ�,�Lf��s�0�$��S��Wqn�ƪ�1I�t=PI�_�/�BJ�_�e٢�^%�I�c��7�0�U\�EE�������/�\$�����$�E+\h
u�c������S��c(�7G3��OZy��[�}ti(Ij�5�v/�u��Ft+�߼NZ�ص���O���|Ր�Gs�>�����j�?�C���������[�gs�u���w�p�d%����YR�Ov�2�#��]��{��(�h��sf��@]z�o��W�8�U��E��z[��r�vd�e�@�0E�O�
���p�w�k�l��e��%,�����]`��������ȗAZ���N�T7#�GW�=K�~�N$�0u��d���6"r����-bg��q���u&���.����L����k/`�
7Q͚����l4[ t�ꌵ��|����/h����;x�/c\xR@��>(d,���,c j�~_/��I�n��a���S<ds>A�Hچk���)"T)6RȖ��߭����$���>��j���
��%v������)��E����S���S����A ��(
% ��5A��8z���C���,�7u��F㎮!&��������B��nBZrd��I���-���,��Go� ��9�U-�Zٛ�}Yz �Et&��WON�����*i_�ʻ&,U�CC����JH����ƾS3�o@ؗ�C�!GrX&��$#�K��rD�Z�Dw)�6�}��L�)����3~L3V�Y� �N��Z� iDA���lc�O��'M!��^�0lN��F��}��X(��3�0���9�kށ�����I��<���ƹ�3B������9^ �	5��wɸ�I4�U��M�%�}GpP�b�s$%�C��ϮfG�g'|˙ �����`�M1����֦�B2<F"����3%��JDQ7�����x��W8�_��%�B
�d�;��H���c�L8];�=� -i]��`0է4�E�FL}�>d;��-%����ʙS�܀��Z��I ��ҿi#$'��q����ؔyo��H����@~�k�0����ʯ�~X� �,.�]J��eJ�������w ����B�������Q6ᘱ�q��PK�&�
�ؗc�����;��qf�'��a\�{�XRD���zҦ�����9�S*��]-~�nֆ�X�ېVb�s�.�B�/��2CcH�ȿW Vf���D��T�'?Q��I�706RY��W��@��u��i�d�3[n�S6.���WػO�ǹ�0�z�5��	2���֒�o��j� �� C
�E�G���V�h����m]N���>�s��@&Wmd��sa�ʘ�<��r+��qK��5W<���`'��M�V���&�n�@d?�(�y��A�n�Xb�_�v�DQ��(ZLG�eeR��_X��u{�U%���V�����~hg��r�{�j�L�G��D��$�|�\�y�� �����!6`Ws H�dReߣ����;�td�a�%�Oބ7���p�[��q]��is�v�ݰŷ7��3F|�/<#��Yu����7��-���"]P��ku|����{X��T%�x0����r�� �5聕��oEf�Y�.T�<ބ����Z�r�R[�B�c|�&X�:������8ď��}e���� u5B�Bu�F}xJ�t��l*�P����[� �!��Ci5B��Y]��>�{�������( �IX"�n�$��bC��
Y��|H��\�2�dM���xj(���(%5��� F��$sJ�d��v���tm��33���T0�'�F��>G����8���Zӷ឴l]����G֥�SM�H\B݈T2��c�\�)���]F�����	�
g)�c��Z*Y�Q�ʴ�WӱP4�|Y�u�i	{�y�ǽ���/Tq� f��y���g߉����9�Z���tD��A�Nm��cm�� ���è/=��>��kɑ����[j�m���<!�u��	V�ƺ)��(���*Qe2�`&��&���������j]
�r&2�˄����+b����Ϡ��g�$��e!Ǫ� X�~�l�e��������5����U����jzvE�2��$L"٭�Qv��`2C��Zf>|Y�J�%�P���_(r����۩��=2x�;:��b�8�[5S�������pu8�c0l�N��r��Ho��s���1����ą��=��1Ļ�\?��/c�̯�l�8o(Z��F��Q/��v���/W�ӌ)Ux���|���h���^�ͺ�^���,�k/j���bj$�uF9�Q7N�|�����}c�Ҩy
|��	vߒ��/��[�����a�#�3�ē���ba���GvM��������q�[\��[��ڧ��xZ*�(d�@�1�w��`7���EjO�垍���[ہžS�6���B\$�0Fz�����R�[�����O�`Y�AZ��X.�qUeZ�Q�E��M��[�h����p��,�������K����-�K

�x��'�	����ײY�=hE|�yG��ǵ��`>�g��SW<�������y�W),�K*��P���c��}�.F�thJ��y�6�#ExTe!=���HB�l�䆓'��j�b�\!��։���
D�(����Uev���۳���j{o�$��⢲S�����h�,�Ʒn�����:�T���Bm-�L�(RB����Q�/��7��U,�Q+]�U�M��
���V%_UͤF�����hB��kƒ%�q�8�ƪ�N�fY�߳%H.Y��Z���BDIS����k�s<?@�x�5,
�1eL�r{�_��t���fh����I��hʄى�B�L��4��Q!l�Oږ��
��`x�~~�q���=L��"���0�����D
y("�TvZ�x��GT榘����I�������Kp���V���M���G6Z2�W�t0�?f�*�f1�U�7O�y����ur\��u!����]�(̳T �Z��uh�i�D�v�Cd�����K����'���y��h�X����y��P�z����r�b�'YQ4�����Yd��2��8��W����D^�$Jxu���%n��6�Vy�˜�P�"u�ӧ������Q�Be`��/�����2���gI5�J�}����o�� ���2�\1�T��9��:ibQ�m.�k��Em3��+�޷�
�AI�&��=�QO�Z���n).[�C1�.���������v��]���
�y���!�&趷z�������A�"��4&���3}����^P���[l�İ�XL�F=�M��w���}�H�(����*u�Fp1j_�C:c�7��������&Lҁi.ܠ��������o=7��4�.�OFڠ�M�YDj=슎���bΧB�/�H��'����cs��d�N�B�Ǐۤ��$��!N���z{h�� 0�_0��k���:��Rh�!ې�^?�pR�k������I}������W� 6}kU⯳���*�Ȇ�]�晡z����Yo�-��p}�W������o��/u",��Mv�pPE��zwrmP|�k��:#Sx���3j�}Ħ�D:�0�� ݒ�,�M�wF�7M��m*%a�)���S�����C[�I)��Og��d��-\�/.����F}��m8�4k���2�A��-���"zZX����*I�o~E��r�)b=M.�\]&���P�7��M�p�9p�ֆ�ưZ=�'��q��ٟ]�hK>�/�PH���=I3)b������bQ���K+iS05�?~ąz�钥�	5t8�5%]@�)�kca�e�S�@3o�t�����zZ�:���H^#�=�M	���,t��}�������#kWע�&ME�dj�6�\��P�(-���]�x.+1��*z��k��H
���W�jy�`2YfN?���-����N5�4�d*������"��\0������?K���g��~G�3�)h����/�&(Nd�Ǥ�2���0ܟ���#_�~�ˀ�1��7k��D���
1�ub�+J* ��R�t�����а'>�{H�#��� �Z��j|v��u=�e%�}O�C��Z>V�NF�G��o	�}���%TED�մoC`�AС�h+��E2I�kT����qږ��������=���V��T�yR�R���r�@���b뼒k���'��C�J�ʠ��֦���ș��'��H�X%�m��;#�Bj���O��U'~2�]���!k<A���IS±�~��Eg�@�_�f����(��%��W'� 3�nI&�ތ���#�}��k�mW���cj�k����	#{�Z_�u|8t�b��wF_,��]�v�L�ċ���v����CZ�챻{FhO�Ό|�P�U3��~+�[r*���0ݭ�A̺9�GT{nη��k}��O��I�!lt��f��g�)��a� [�9�p4~�O�W7�"L�п11@�F4߻B+>�	�d��#;�Ar@'�cA��Sf�2ʐF結��4�ط��/CIaӁ-�K�8�S���ǆ�B�a�rg����a����\�,�"����=�1׉���[�}S|MGqB�U�r�u�f��/
�9��9=ɛew2��V��u�!��˛9F�hR}k���)P�$��'E�,�#s�ˎ�S��^H��(!��W�J�׋� 	�^���u�'��/X,M.^K���uᱽ�t������\�Z�ke]�n,��^��-�o� ��K������r�����#Ֆ���RR{D����˔�f}��=��.;�ǣ�0)��e�Y��g�)�]�;Y�xngNĵ�rA�_�9�5��P�O�^�fܒx�]���x��������h�@[�#��y��������6[��v�����	��J���/��̗N�@+�Y�Z��5ۂIEm|K��o ?l4��|�#*$�Ѐ:���TXLJ@a�(��&���]�5W#L<��b*A��
�����/1�90�~��1a�T�K�w�������H�C�'Iz!%)r�J���{>�R?ӕ�;JƬ#⌱���5�]0w�nM��7K<W$���EIV�Ȭ����|h��ϢN��B.��E��hA��f	;<ޓ �I�-�pz��?sdȓ�r(3`���������И�^�?����	/fI����z��ؤ�*�'-I��R2[��T����ڕ��+��<�Y]��v��1����b� (�G2�Р����y�;eل^��i��u2(�q�-�0-s0p�y��աޡ[�jC߶g�4�Z<�4*�b!�	�$B�#�ا����lC&,�B���*�x�| ��G�l)�˄M�دg#ѕl(��K�@�"<��&��$6��9��J�ײ�E ���h"KJ1I����5=A���P���ּ'��>��ѵ�@žߠ@'���(�L�y�բ�[����j���W�B�W6�@<\iӤSU8� �nC9�}��:���u�	R��08�]n�|���񐟅D0�m�K�{�oxދa��kƖ�?��83���*�$U��l�p��ڂ0��h�"Y^��2vz���}67��hq-����8=����Ȏ�T>������%�,j��뛘���Z=�.yH=&j���<�n�wDn��4i�-�i�����%�h0���:�_��ے���Z��Ȗ~�#�����dM���݉���s2͋:�@߀���e�U�?x)��=^"����m�=��k�q-x]�`��Io��Ҳt���K�p���P�WoȊj0�|�Y�RbpeuO&��ېG�����1;����iC��@��o��@��:E�"u�u����ߋl�I�7(�*o����l)�)���pβlMd��.�7S�L���$)���>�5R��~��Aq��^���R�(�n�c�57�5i�Ŭ�e�����y�� �^��9��4%l��tE,�3u+�VX��<�/YO
�搸����>dV�7Ud\̨XO�݌�cn�K�)s
�����
ME�b���T���T]4r'K���y1��u�Q�9�षB�L�\���"l )i�3*�C��u���`Y��R�CI6�n�A��[�ɚ}�7d��T2�J�+$�\xv$�᢮��]�J�D~]����`=$u-.�kMg���MA0������ `���>7�ي>��"��H��D���,���eX�]�$�`�V��R>W�ծ�Ŕ$�X6��)<��
��6��)��ڋ�~'�˫:�|s�Gt���Ig^�`��N�6�	HB#E����5���
-�P)���,�w� ��6���K�%�/������	�w3�Th��y�J!ޡ�$*�A���d�Ngo~�S��S�zm 	���80�=���m������W�c�`g��N���\,�Ѵ��~��Mwyb��vX���ۘ��=;Dt��nd\_�0K%�B�8�S6��N~j���@?���;�&���i{�X,O��s�0k��-�6�
s>���8H�V$}��G��I��rYf�ۺ�uI�us������f�)�^𱣛�\I
\|�T��L������/6͕2��8�����}����}����Tw�{Ԩ������U{��Iʁ��y�3ȉm�d���?8Q ����c��:%�J�K�߾
	�YbxMCnXjČ#�
�sN�w�3{�T%"*�D�-��ʆ->�KVX����yr���Ż���XQߌ����6B��v��$��z�����W�AYxq�T&;�w���!�T���p��
�z�&�f-4������̾0��t ����d�f���U�u/\�8���Thj�Y��~������u�ьDi��޻g�?;�C�0��	/ j�ο-��l�T�U���Q>�������Oѝ��?`Q>zT+n`������"��]�t��2P����%����S��Al B� �c~�;wM��hW��=��}IX<:O��75B�ߪ!���)On��r���F|V\��7��o��۽�"�#���3bY�^1�c���G�e.%ڢF��f����l�y�Sy�Rً:�� ���5�CՂ��^�c��&)λ�<wH�-���r����:�Q-�?<Q�H�O�P�6'Uj�0��G��y3m�zU��c�6v݌'����Y�s�����.�?�������G9��{�U�b���qM�"�<zk���B��`	Q6�V�x��Q��(�ދ]}��b�M�c>Y�3�-3��<RbW�#�m���&� {w�����\������[Ӂ���	�E��+D!��aGq��&w���p�/9|���X�%�}q�`���!P	s[P&�ߎB �4���uEN�6[	U�0����n,i̨+��A����7-��ձs�Qo�s�/k����4�}�s4?��kQ{+��H��`��tA*���>@��ʺ��P<�����RF��/s4Y��(�:���(��v��_X������OEM!��c��=7噽���s�y��~�!��cV/m���<l��}�����k�*�(�czr��pOU�0�N��jS[Mf3YG�:�{P�7O\L��! U>�P?�,&�x�{��J;�iD�7�b���#f~(�(�jȀ;Ig��v�1A%��YJ�:���K�~����K��z�rx��>�%2׃�z��6o��$�7h;Z��:5�v�*;/`;���$�_gN3ۥIj� ��'�G9W-?��2�ʁ^�C�K�M�M�n$Ҡ�_{�G��R-�эot�q ��l<d�'L�#t����z����H�?� x��Nlrxe��|�Vr{o��$生�?���_�cq��8�`���ܡ�h�ёO�l���
�	ym�'�7�2s}:�jV�K5l����j����������ٶ�8%�|;�8�;���@�����$�4�)s#KJlF}/����o�ږ&t�!�C[���6 y�ۻ��y��� �ξX��H`��;��z+	���0k1*[	q����k���C�68Ď���۵�0U�V�Yre9l�G�c�+R;~шW�&���׷�$���GC?SZ���~��Y�g\,��h3��\���/$o�:e�w���C�s�U�B�[o�Cl�h�M��0^'
b�E	c��CT*�Y4�,�%�����r?���Î�<��e��U�0bI~���=i���( )��|8��¸ްgG�h5]u�VUK�<Dbiy {آH&4?�ȹ�X�����1��l�4�g �ۛRG+�b�nn���^0,z�1����>^����a��=A��3�0Wq�X�ͽ�ٹ�k3�W�K44Pt�����3.�����7m�
�Q�j�`�S����*�%:����⁬ь��7Y���'~�?ԳxG,E�Az{����0��L��M���u�S�F�sV�_��l� f�bc����ǋ���v��K�`�l����|��2X��3�J!0L��;,lLvN{Z�!:0e��T9���˥*{~��ʉ;����}���s	蝈�F_
Ȍ��1k��9��|����Z|qj�>���`�3�s ���;�f9��JL�E�܋a}`\͐�g&u��@nҀ?)Z��l55�?��m][B�/�>VΏL����?��z�,�Wn��:*S
� ZWh���[�hR$�@t\<�K��5�z����c�!����e��6 �z��U'Ȍ�-G����H=n�^����S��C����s�Zښ�N������ 9���)plod��y �潖�|���-6��º#�P)v�i�v�]7����{T���L�EÙ^�h9�ef�k[�[�F��s8t)�������2v�-�`8�ֈT��-��yLƌ�'h���Y�C��Nϑ��:���J�u�a�'<��0ZI�7���,U�j�wc��ޜeT,|ɚ	F"����\"J�#M*5��ł� �_g���.G��Ǐ��ŀ{
m �cC�֑�ܡk��ҳd��:�xٱ���9@:jUp�Ɍ$�/vJ\�������Cs�j���J�����ƏHi�����m�,i�j�#���&�������쾣�iT������m�u1J�k<��Y(�p~�E��Z�7�D�N}�h����{̶�^<��1iy�m�}��.��)���}#{r������<��7򕍾b���[�5���ŷd���'h��9����?�C3���
�"f�@ ��ջ�l�B�͸Aj_�cbUi��<=�1�������Z5�ўc��:���t��d�PdS�8*jS�&���Gf�3�N�[���p�> �qi�1���4u�/��0��X�7wN��Z�hK��H����$����qm�+���/�n�A^�E���y͗TXS�Z�4t��Tt]���Ã�����Ɵ��g6��_w�w��]����{�[Ĺ�(�[O�N��ٔ��.Ӏ�  n��r����H���p�x�&�ḍTc�	T�Cn'#^YwW.їn�ڢ�=��s��OL��
a�%�1-b���[�*�v,��(�`.S<R�U/y�,�^N[��
���V�c!�G�����;<�g��K��5�с�_����Do��V_�:��Qc�+/w!�ޥ���%��Nf��g�U�G���9�ݜ��5��58�'�"ޖ���k�u*���۹�Ԟf�;���щd��w�7�j�>�UOlw�k�6h��B�gAĜ�5����&���^�~k�݇f��rK�U���Ta�j�8#Qiȑ��^���д5��_�T���,_g����.�
Ah���ཁ<�Bf;���#1f�m�fjA/@֊��o�e��� }�o�ٕ`/�(@Z n��p��:T� 0�p�^=P�H���CA��I�޿Z&��NM�a��d$1E�����}]_�a�݂��\�vU;z��[J����(�I�ƌi'B[:/��@�)D:�{^%x�΀�@32EJ:���lh�}.S.�����r-�w"ԋ_ߜ�o��p 0�:)T�!S��O���^�J���R�n;����� ��� -	�N���`��Zdy{��{��C��N� �������-`K_&)I)���ȁ���N�o�{�?�ͥ�EZKf�Ad{�T#d�R�q?��d7���÷���EJ$�/����4��E��Lz�a�n1���04��������M��	N}���fE̮��e/���8hW�]�<�G�n���׌����sC��;������Я���h\��jxOZ�}��� �>��e{���*�tb;{b��|{�n�&�J��i�s���`~�!p6L�wF�����B_��&իY�]�C����5���"����߾�$����SxU���,ꃼ�p߇����Mz�j��:��Pt��	w[�B�$זJ��`�t9~V&��y��cO���4��K)�|�~���5��6��Ruh����**\��x�Չ4���>��n'*�,b���6C3?|�
K���pI�3�(��6e�0�!iP?y�\�[��v�����zu٣�+6���r4��P8)&#�xH_X(3���[���b�Ys$�{"Ɗ�ǘ��{$�����35?�cXK�0Z
v���ǰ�ojː=��*��_�i4�.w�jm�x�����O�dH�h��:� ?[�ړ|0����Z��[�;+��i��sJbg9��ц�w��#4��f�U�_������Ae���4H^}
|M[3�ݛ�Y6�����40Բ�(�i�Tq�a'K��BUz�=ok�T�hm�F8���w^N;Uŭ�_��%���f��$��Y@�9R������������ʼ�E���a#=���:a2���5�!����f}��n����C�x��N�7�y_�cQАi�h��a�N'ƌ�D���&W��zc�e��D��M���7h(J��gC~��,�oJd<�î9Ր䛻����C��~9I����VX1`#���5��0B���#�2�=F K�k��O;��V�=�\���p��=�����Fߥ���\ �>��|x�oٮ|��g0^���	�Ë4c��P�8�������yxly�b#�����"Y%��r��h"��b�!(���JF3S�J����Bs2�ɤ4�h����*�hq�Z���D��s�Y��-�b�AY�d�k�s���m��E0�+d�t���C�*-�j���7�r��ɡ��I���>8B��9�w��Jj�}�-�HkR��e�)��S����C3?7p-H!zXkf֋br��԰����l'wl:���P�W�;�8�3�>�J�\*m��y�5��a��E������h��_�VM���|r~����%��M�D�$,�/di_��<�a��S�M%��������a/�
Q
l9x�)��{:uzo��NKccZPʣ���)x��<mؑ�:�j���ڞ+I�π���P-�Z��ЗBU�'�����A��jn2z�TY���*�����Ԍ���oj��6o��.�N�+��e94|1�~oڽC���.�R)F�~D�D۩�W{� Ϡ�$�95i��������������]X�p^���Ů��%F z`�s:�)�����7��Y��� ��AۿJs��E7p'����je5��ݭ�ݕvLL�_��v��2��ҽ�f�v�hVfƺ��*R�b���ź����')�OL3����!����{\")��2#F�~`�b@4}�A?�OĂ��=Q#�����Ϣե��{�Ȳ��+��� ��P��\�la���c�+t �� ��-�>��lRn�4�Z�}��ӊѦJ�KO�����:3q���!#�@�U������A�9�ickd� ����"72��㵤��}�uCэ~�ÿ�)���#�ٟ��g{�so����g��C/��؃	{�;�!�["���؄�c��3�"�Y���8�H�ko6=�.�	~��+@F��V�+�c7��זސyI���;M�B�n<ɑ���8�kC>�IF��<4�sr��9�EmNT�K-_ρ��oJі��y2���TV�v9$4���2:KM�3� Pz�Z=-�C�V"�O�����r�_��A��lc`��ʓ�4z�JGnAb�S�^X�n��ݧ[�B6��%���	S4\��{��7L���[pLt[	�� B�R��;�jE�M�u�`*p���m�Y�t�TE^nϖ�6軭����L�Fv��,�.��z��w���ˉ"C�HW�#K�	��G"�
i��6��t�-%Kǳ�ِ
�}���[u��}��z
h��G ���鼥n�
��TX%0�	�q���*$|PI(��8P�,���%;����s�o���R��*[�'C�*ViG�����z6�ei�Z�qH'z2���B���o"B��z��g:����)H|[�A#72����Nts����zC;!�5V�����j���8������:����bw��9�z,J��֏r�{)4���O��B9�
�\�.4�=�>sI��*��-n>h�u��֚x��xC{�GW�����0[�d>��j=fKG~�/��C��3Z��p'�n��FG�����Ɋ�є�<��@����>���ǐ	�1fG)�r�u
� �2�#��~@	kzZ� ���PW� �7�^a�Е &1���\�V`���B�iA]�W `��^ɧ�0�h�L�k.>[O,=gI��@8W��U��u�s�g���(sp����[TMu*ݎ6�to�-�b���(�-@�;��hCv�Ia}[�֩-&�
�j*x(=I��al]&�(9]�Ե<gh�v��H*�x�Ikv�i��Ƕ�G� ��3����{�X��t���P��~��c��ܥ^�b���AɹA#R̤�dK���1:j���R����Tj���J��E(0�_Z�8��I�p����.4�QXohT�lᑿ�\�޷���3bOPV(Frz�FH�� :����?q�zVE!&ՠ#��B�sQ�O�yB�4d�Ǒ����Cz�P�l��D k�~UJKߛz�.ݩE���t�|6�����*r4�5&u+�<�ۚp�1���5����^'!8W#8�y�OĶ�R��	J�B�ρٮ���Xi���;"z��j��V"5�T�|���+&���m�x�C�G>���V��~跖��h�@�)�^_+RT�����2��7T����d���{Z�De��b�0�θ�I˝�'�Ƌ��#t;�9�4@{s��52s���b$��l� 8bU[$��j��p.Ϧ��0փt�CF��0J
�9YF䋿��r�kr�`�{h.��,���:j��A��3�����O������t�z��[7(w���Rwb���&]1ь�z����s�>��I��h�:ծ&�c�کZ�9{PB�S#ԡv�h��|٬3�x� � �H�|
�y /O)@S������:O��J�M�F�~���-�S+V�^ul��E�`9^��[��y�WP@�}�~�Z��1��P߯X�J��}\/�z(���V׬!lXG�`!���y���4�f�R��ZU�K�z2�՜�b��a�mwp�v����h��`��k/�;&�N����C�ռ꬟ĚC
��|CH*0I%|�z`���n|��Q,�U�{��k�V����R�
C�ϑ���T������?���F|��]@�4R��Da��F3���̿��	�,G|#���DE
�;�R)V:��.�g�3f>�B�lV�5_N6+?�2���}��Wq*�|�����!	��ڗ`��~��C	�v�޾
�停lV�]cP�:Gk�D��r ��E�iD'��ꛉ��nl����I�����n��vV�`�W�.�(���`_xg$���f��˅�߀�`M���ax}���)��cI�n���7��#��{��%=J�f@Ϸ�L��X֬���4|�~p�^���2�h�r���
ߕ����q..�-ԓ�F�{��4,��w!c��r��<^"�_YE����|�N6ź*
�&'PԀ�]�� XS�nxT���!q��<\�M4!���nq=�*�Դ��WS�6��3�}����
��c��@kn�(��,�	��kI��ħbH��;��W�ٵADAŞ�k`���O�X}�w
<����HE:.����@&E�dt�A���M�b�kQ���^X�͹˩� ��L��m/�}��l�w
�n?�$�|�m1�te�B���ٱ;"�	�N��-�u���$��lQ����˦��(r*]r�o��O�ۦ�S<8o�s��습�$wr�v"���a����6���FD\��Y)(D�gg���lm�r����Ͻ��h;���w�]R}8��O���Hw�H�Q��mS:�Z�����.������%^3��h��؃��2���<T��F�槫�P]�����?��9\�n����i�Zih�g#WD 2�Rs���t�ଷ����%e��6%��c�K��P��o����C�B-�[�W�0�ӕE��1!�Ѳ�D��η����a��^�gE���a�2�
<�(��l��5N|چ��s#�*M��n1`����صwe�Q$���!�[�<b~�W�<N��?v=�E�J�=�J��� ~3e���J^AQ�=;�j��S�A�A��o��e8��
��L������5�\W	�-��J獉x��Y'���=6}�Y{�������28���a$���|��j��5��1ٰ��~�'�tpg��J>����b���o`ޒ~-~�u��n��ﵧ���RAjW~e�����֘�9�����-�B9J�7_��D#�yG��S�߸��m[ݘ��/0+}2}�]����k��]��I�!�����/���L�%!@s,�����
�\���-c\Z_(�����?��E���uH���$ ֢�� (*��n��đ���󕫑R��_�S�:��7�<Ei�Ɲ�{�Tt�Xh^J��^o�C�z��°8Ek4���"ɖ�'K`/��XJt����� \����̇�Oq��3�3$"O�i=�.�i��z�(, w�KA�S-�
{E�#3)��W�:71�}�ǂ���R�@��.�?�wb�K0l����3��O<Wn��g[I �:Ga-nk��D�x�+�
x�Îw���b��@=��C���`N��)���vB�(i"�s`�����2��71�%Xo��Ȳre#1��{OuFV"��ظ \X�qZ�
�Z���7'4T������\�����G`�Q�L&0�[b�fx�fZ������݈�e�GO��m.i�Ț����D�*Ȯ����h�z�����i�/�qL�hp�w�l���@'�o���}�����:Uc�"��ݍ9[�ǻs1eTZ���(�EU`~l:���7���'"z��CyQ=�����* � *��0�q���N����r�:m���YƢ���?��u�r73iJ�{~�xҌ�;7L��)�B�.N$�.��-P����Y�o��W��)w���U���|A݋�
��>v�A�\���a��t9
�]�2S��0*t�q��aӷ7���|��^LA���Lg^j������Q�_�B�㑲����+Q�P;K���ߟ��Z�H��iGŚ���Qςh~I�=��5�O��Ů��V���������r�]T��䪻�T��ؒ�Uzqr\u��-}"�ߢ�(d,"�P��7���b�J�yC!��<z;:
�=�2��R*hsiY8 b�Z�
kR��y�jKg�H���R���CZ|"���(U�q���3s\u��<��q���au%�nHQ�/(V��T��ړ�g�_��$v���M��l���c;��p�`R��ڡ!�4�e�<;�B"���m�v��M�:�s� t��!e2��F�s���r���Ȯ[I��R����5^v!�^�|��U�SG/�D\��	
��VZ���|>�Q��8��/$�����Ơ?�H�,ڞ����8#�3�h=j�:�K�[�C/Z-a�@RjJS�����k��6aX��I��q[Q��x*}���g�@y�2E���3�<��r������	K���8����� ��kS{�8�{�B �F��\��^�)�%�KevB���*ǆ1e*�zv�]�
o>0�A`(��y'��G�f�&�����{�@�M���~N5D�����q	[|¨,*��<K+B�K��FޔJ(8\=/�^�]'_��`܏-N�*���A�oZ�c1E���H)~���,��KLeL�#gnF4y�BLq�#��s�u�#[�������r�����B�T��F0zЃf�_��L՜��f:\���@���3�=8v�]Q�ѸOi�F#�4>/Mڵ�*ǄK�����tiZ���ZS`��w�z~l���ݺ%��z���}�s6�j:��7'�|.�D��nQ�ْAlLM�R������S�N�/�ٮ^X���ߡKb?2 ��[dq�F�:�b5�����NW~��z�7A�bW��U\b�K �.i�#�tSq�&L"i�ѽ=y�'��f�&d}*�� v-���WQ�⹂ɥц���qR�8������@&�GH�� V�!���BÌ�xK���|��l�^���I���3M���Z�)x�w��U���QE^�L��}uw�<d����)|���WG��k�F�1�%�(�own���Uk}�~Q�i�2$[EKd�m$�\�Y�@���32>�`��g����_�t��Z�E�.<�Q���3�q��J�%k�َd����ى�d���L ;U���5D
$M���D�3�3�뿥%��"���!�^8t��1m�
��!����"�S]W�lit���ck�Q����߉մ�bnF`r9�5s���\����ĽE�8�G1��Í�s7�9��+����1v���a���Þ^ZX�h��]�*}@u�>���@B�nَ@����_tG�µ�|?kK���$��,T�6GϪ���}l�w6�
sz5^I�G8�M�!�.
����]��~�زkȟ�L�Z�cbhJ��FsXO��s4.��Zt
�����opɢ�J�cE�#!��qq�)�Ii�ڢ1�)m�U�[��P��&���.��+��/'���įzj�Y_�$a]&��T����`!,p����&	�q�`S#���n_e�1��s8.q���4����n�����9÷+xHMuI��a*d��Q7sAH�J���[CK�,�q�Y�>�"�D��i�B��m�Jb,B�$��^�9���c���W-��$6'O����_��dr� Ho�v�7�CR��rt<$��>�����fN���Sdx=�!�0�� uk�pp=%y�R��@i��$��3���Z\����@m#��4���U�+�q1A�p�Lz�­=���p�V����ANQ�����p�ڹ��Q8U,w�0���/SA�� �����>F�Yk��pE��%vR���� ��s]�cǒ��F(��KЪ��uO���p�� ���o�8��j��H���X?�M��q���/�9���Iu��j��!D1�L�m*O��ɘF6K������iG���
��R������(ο������'�7w�^��\2�)^�+�nIE}lZK@\�F��BQ�.��4d�{�BKd��YȄ�+�w���	ԁm�
�S��z�\6��#���u'�(o�Vy�f��i�TB�ߥ��Q�f(vCzaͤ�,���iS�X��M�&�קM�A�3Ok4�ן�3��X0�Q���}
M��ߜww�֢�����0�-�y�EΔB���������a�!����d�p�^]	E�;�9����
��.���f��0{e���(�1G�7)@⛈����斻�d��l��*���zX@D��
\b�S�
C�u�}���9?��.�mW��f�v7(9�,q>n��W]��ٟ���]�<c�~g�7B��V�m3��+V[����"
��]�:���5PѢ�ȷ �^�pU,�5g���r��->:��HA]���l�C���S�ԥ�,��>����>+�}�Ǻ0��z@#����ᨨ[%�֥:��W�����H֚`yVE/�jϘ��9'!�ΓѦ���y�̢�����:�RM�[�����e!�^�
�eT*��-�i���J}L5��ǋ�'���Q~KD����1Sul����e�؟�>�8� S��}�i[���YuVO!��q�lP%>��X& ,�eխ�S��媶SC���'��+�+'5�YAf�Y2����k�t8i}��h��Ț�cp"8b�'����+�!q�#
�t*�K��S�_g�@�W.|�>,O�1��>���^stJ�Q�{�px߄s'zNW嘝���"�G��Pq�p��L�&&��lݝ_�!]0�c���#�MWf�o��:2��� F���aL���S�QZ����K[���d�Qq�P�a�)���k%��ޞ��$g/�[*�#��	�g�^� ��������(�y`:�:V�����k@�b@ :����s�ěo�#Y~7��!�l��s'������z��3
@Y?G�Q�������W�z��U(����/i6�dCy+b��ӣ#�6�V'���P�-V;�+�`k�%�"x� �S��.��ٜ93�Tj�`O��yR>��UV�=��Mӱ���?^Z�}#�Cj� ߈e�v��[�]��$ǖ񄐌�
�.j�JlA��EY�F4L�ω֫��=� t��K��S�n8�q����j�K��k�&� ��>�6
��	���H��o�\la;��0�X���qO�q�@���:�����}<Z�ڴ*���g��=��R�H�AQO��jX�S ��5z*��R`i��GIR�����MF����gg�E*Ҧ���d��	*��BC����4M,.x#�jP���~@������$Z��������[(�߀�|=p`�&&���KM��^���ހ���lmG�TO���R���]�6�4�mD?��$q�X�s�d���i 6��C%��}(X�	��]�!}��Z�;�9u=���)�a�����$ f1���^�����O��;v~���9a�Maev���s�E	$FS����|�Tܖ�,e�,��`��H�����J�=��y<\g��K� �nQK��6��'���
٫yF��}�[����h��I�U�FsgC����jL��䶰�>"eD�ZJ�lT��߁I�ۺ�2]��u ���(�48�L4���pu���[f#����3��d��4����򀴵�6�1�����2�	�vi_Us�
/m:�(՟N^����/��$�� �j��7�7�DF�R�_� y�UZ�����j��j.{��H�Wr�NT�)�ϹI���K@x�h�Y�f�B���4�������qS�-oo�a�(6V7�_�ϸ9���G��|
�z����,�X����&�.��CLA@��"z
ӊ�j7��� f�N��F�!u�/Q�LF�D�K����פ!J����_x����k��J�T�xfd!����y�����;ԻÛ�
w��<��]H�,�<��B|/Zg�dN�[�tUp���������IR��9f ꯓ�x8��Llد�Ӊ�4���a�{<�+��{����
�\4�Xдz�#�B*���E:h�x����f�bZ��@�
�H��Cٲ��5w�\L���u��w��>�6
�q�J?#��Z����%��@غ��g���6A��Cwy�Sh�wK�.��v8����Bn�k1�ݱit�-�y���!*�Ļh2	�;~2)����錥�}.\.��TT��?@U��C��3aA�>)��V'i�M�T
__�}�Ж�'�rI��(��M#�h��gf������>��Co�t$��~Z�P�3�jUS�g+%8�������1���֯2��s�9���5�j/J�Ι)q#�������4U��Xj��x�I�TPB"�!����_/���Qsb��>X�����y���⑇�4����<���	�?41�����u������R��	T!(<���6��K��o��wx�Y9��3��YqN���Bٯޱ�����f�.,�j�����B�ad\�4��vu�q�"�`}�dF����;!�� �\��$��~�9Ƀ��Q��ȸj�a�`6�Z��E�qЮBAMr�{��_i%�/�r����Lԩ^�Q����n��~���G�e}gW��1EY{�jU7�@��%�-l��d�AQ%�[�,�՛�U�5�z���+��9ɓ���ӗr=�,�KW\Hs��W8�@��l�,Q	�!h�BR����_�D�ع{�Mq�[�@��Մ;Rд렺A��"�A��Ŭ]��?��:�n:�h��1�����!�� cF�C��	{�����+H�ȳ+��#e�n����/!��
p��\�DFc�|I�#���Z����p)GW���@���J���\;u�rlĬ�-饄��@����FbưXu2����`I�u����o*%,bW�Kl��S�!����q<v1�B���+��y�*q��O O��i�iiK��5X��A�F5Z�թ<�Z��0���wL,bخ���.$w[{!�#����}��ά�@?N���7�X��`���
_�a���=&rs��;_@��i�bĥ�����9Ul��y(̣�q��0~��2��]}�^�Rde��.�
n�߸��'���@�;�q�%�UO�=q0j�u�%g)�� :#�#�`�rM`6&q���}�YQ�.��)���V��� ���ݿƨ�?����K2�_�ݿ���s�}��e��gP1��R��!-̄�h��X�e���{���恈rU_]I]��7IrƠr�&*�e6���f�7J��qWQc�!�;�	a��[�WJ�,��tR=c>J-�&��0�pu��C�5'�xgn��Wk��ΈuƂ�\�IE/�w�M�J�8Rt�˿	��'���N�<!���7�Ǆ L�ds[������N��S�n3�ȯ���}�����z�I���PY�(t��'JD�8�&&�Tt�o���r������/���N!��	Cj����p��(.�+�3������]��
c�$i�@�j/���� ��.W�f��C��m��Mfu؄s�Q�z3��c^�94��Hi����2U�!p�M��@F�@�6ιL�j9��K����q�Rn��r7;�j�_c/�\�$��i��M�c��S�b�0y����:�Y����InYl"O��4sC�����6�65wg��^N6��Qia���Z��R���?q���ڦ/љ��>V�x�GL��6bJ*o�N���Wk��+�t?ɉ����AE�gߦ�gok#�=�c3
n?n҈������e�y&���&�f��|绿�z��f�!�D��<��?�bR;'^�E�|.��������v�� )����y�ז�c��ko�a��T+_�#J:�?�a!n:f�|Pu4ñi�DJt�!-�Q&�,�Xp��8����:D�S̞�c�Y������!�Z>A�օә� �f-�F�KΟ�Y�j�Wh3�P��̷��.�6A�s�o��H���%9X�;*ﾬA;v��:9b�C.�*�!>~Ox���3����Z�s���s��_��đ�~ ��P�Oa���uGY T:
Kdg{��΂���4�٨9O�K��4�߁���Y�>H��͛th����M��iz$��X�7��E�а`�W��<���gw�=��k��}E����+�`�7pk����Օ�9@,��`��B����n���J�`�l�H
f��4�W3�z��ƭ
�ó� �Y��o�,X-�5N8K��� ���:|`x�y����Ck�j4���w���*(��)�,�5F(��-��1�+cYOrkUfp���}�����7����^��N�үVa����u��Ôx=��F���*,W�N���l
����3|�S����u�5�Ѻ�d�8)u��ޒΖ+��ޫm&sq�w|�����[�C;��͝_�����8^S�
Ilx(��{��+U�>���1|x�@h�a�Q>I�I/^��jE/|��}y�	�,�֯���~ؚ�ؠ9�� 
���f��*�s������4�gʇ�6�)�:\!;�-$�{�;��0�ןW�Zv%��_9���.ĉ�l�l��	��[����rTq��E�~� ��,�\�x@�A���~��.1��PR�
,Vcf����>���m3 6X������3r=lH9��"��3�7:��K'g1�D��a;������yWW��u:���Iؓ,���erЌ��(�{�p���r��ڦ�{/�k�;��s��CE�Z��,[��89�5Xs�a�W���Mx���❠Q�21��,�+]�~�D��rS2/�ϙ����2x`.�wr�vT�xʟ�,��N���4�؍v�L	��51�i�����Cr�����mb�I�dߠ}���i��p/4�/�j?���҉rkĺ�Y�{W���
�1�N<\H*�@�)o*�Є���75����/*�t�OBS�9p� ca=��M	^��ƿƩ���]�b�4�s
�S_�\���uMf�1W�=�vF�)ǻW�P�&u�w@�"Gj��qiՉK��4���M��u,A1޷�6��o�Ŧ߫��ʑ~o��~	����n���gw�P�����<5��IM@t��>.T�]㗡��xa��Ȝp�,�j;esL駈�Ǹ�v"�W��������i&D\��3v.�f)������{��4G�R޾��x���Ov!L�������TI�&�Ƶ8c����V?�W!6+����]�_��"3��Ծ�Q�K��s\�6����gm��0�X��Ii/�B5�u��N���dWg�j�}�.��HW���D�`����,\-�V^���ߠ#)�L��<-u8�Ja͆	�x(����Q.`�`�����/)�w挚S?�4�S)>TC���s�bH�zC�<��J��)ȡ���9	��z�����b�35���_�[�����\������h�a|���G��/�f�-���`.�{�N(�k).�a�?�To�B�6��|�r���Wo��-��x�1?�-�F��D�$F��6L��ؔ��~c T�ߐ2��?t	"����*l1,�����	Sy�&Q�2`dr/�g�������[�h�4bblN�leY��1Oc#?�D�4	P�j�y���]uo!8�z!�ueUE�y Ȋ}�)Ii6Q���νB�D���B8 ֬��[��cǈu�w0��z�G�z_�tV����r���,��v�r�µ!�͝���ׇn�z� RȞ�eL�1�F�P�sfX(��=̷ܥ���J�et��ٯ���J;����U�	�=9**���4?��_�rR��ET2��ԧW�7]�A�-�j���[Cй�^Vt�(k�;,��:
{Ė.�-���?"*WbĒ�=�-AD(� (ȏ��!w�/�wUg�N��M���`E�)bN��c��L�QJ�D"��/m�M0���$��)��wS-xm��_ƻ� ���e��Zω���R�3x⼭���قZ��70a��_s!��'*H�IOI��}f�ҝ�ɫ�돠�s�U��u�μ���P�5�;�c�7UV]���^$��u�~��#���V�p|I@RZ��#�9�>���cxO_�nă��A_ f��������ZK���h�yE�2���T�	��C'�4���%�#�[`��SXV��b!���K��A�������F%����T=�;��v2�\�0m:�Տ���# j��@����;�\�g�g�� M:�E��KC����~"�A˄�%D1ɺ���S�����cm��b�ՠ�ܸ?叜����Yz�C�a�K��$�T��h95B&�h���ix����mB����{��`�T1���'�������;b	xgJ ;Sx;���v6�C]�أ$skm&T���@�����X�<~������Mb�O�;i��*|틯1��U�*���}Fe���Z	��*�c�).o��2}��\�tT�l�y�1н��d����TQ�6��;��]R9��it>d3���C�pvD��O���{�H���!� u�O��u]Ԏ0��6qE@q���!9��82Q�&(��[M~�������K��h�O�=8� 
"�h��p�j��H�k�gG�>�h����"���)����P%`K9U�[�5>����+b�����c<d�'�!b��}��X$�Åm��P*A}V��)[|�l��xwA�Z��0m�Z���@���2&+�;��U�J��N3��&���;t͊��:+�_�"�)rryd5X�( a	����NT��w�����9"�~��?��xW9}57��{B��'�r�|E�U�)t�ߞD@R,>*�B7�bXls�V0��#{tK�o[�]��sl�w�bhR~tLy�����*I�elK���	�Tq��t��,/N󂞵�E��i���O��s��9�wv�OO����6t��CN^2�I��v5�i^�u���W�4�}�iw��X�AU�ߤ��gNB�8�����#~��G=�gi���9lz7�z�V]n�����;L1D�.�f>�H��@q6q,W������BՃ��E)y}���a�f�+�S��ez#Jw�L�d�8c:,[L�\-�&�愇���Z��y
׏I˺}�-=���p�j(���R�v�1�X���0b�޲]i�y�"��{&�h�v�߅���T9FoW١�Y��͹-�fQ�}0k�Ӝ|��%��z�(��}�/:�X�}wM�O^�g)�gh����H�����r���D�֟�K�EW�5����<���J4�/�L=Rp��.n��^�5	�uF� 
��Xh�d�JkN�nI��ć�8#Y�#��pƷ��w�q�cN:s�r
H1h?�t��4Z\�h�~Jn�
�hՍL/�Ww��l�@wp�
��$�Sg����`�Ӽ�x�ɠ�L"l˦\�`��А^�=��ґ�t�t\�q�+�5D~.i������,��l$in�U;�?�}��7����pV�=-�k20Y�w_�Bɱ��������)�t��[�%�[3�H��լ�w��%Gů.�����/��>C����7V|u6��6[9��p%�z���VEǾ&���7��PF���QO�Q{n�6p ���'|��K\�	Pl3	8%��ܺ'�-Z����G!I.���r��o���w1CYWB�&��!�9X.���? ,��ƅw&��[�Cك�G�ݺ� �^=���+���`�!�B�n䌣59h7,�#SrZH�h'�����cpA4���E�F�f���,�&���'�"�{��7q�ǷJ���;Oab�p����������;�9�ִLxnOϋ�q嶤���q��T9�W�%���2�����a�|wL�N��(��FRFSH_Ĝ!�dx�p>%��!�������w���%7"�L#��_�[
3Bɥ����%���Q&N<Q$�����;�1@��d0�6 >R��J��x�gRt�S&�'�����[�\�b#z�4Ž ,f�w�|����ֆnb�M�S:,������ŎE����~����bo7��u��GT��	b�԰F
-ӓ�=A_���G�0�3�Qæ��d��9��	/��|d�QO�� m���y%y��Zgڡ�	�b�p,r/D4��~�0�D�Lz;9'��n%�hf��2식���Ct�W
�ɘ���vߤز��܆��dX���RLV�{S`BG��7/�~0 r��=*o�i���rf�[��=��i�)�w�H�pW$�ܵ>���´�>�-�
(�2�o2�ފn�
&���wGi�J·3۴Lj��Qz�fj����5\�.��H�m�%.���$���#N{Bf���t���wp;��L��o�j���<A5�:�s��O�E	@3��� ']�9Oι�3���8�d�������{��1!7���<���'�&�օ�Y�:i�g���K���A����c�u�N���1��{�=QpkQ�L���pXZ�����fT�=�;�4��}�.1<G��4!K�
�l,����Ru����ЅWBRf�S;']ç|�oX�}*|��1�T��UHq�jmFm���hy$G(hɌm�����?����W$Y*�w���a���u5l��֑�z}{��L����k۶���cU(Q���v]a��8�j�(�/��?|K�W*�`�v�4��*��S}[5K�&�J�YH'״G��M�^��2�Xk����@���h
3��P�2Y6�|Bq�iJ�]z��v�f��[Üj"&2Z��u�.u8SDY$$a���JrPQ,&wJ��$�B��X��[��S]ǫ�Wpe�9�n���?��̍j��T�UM����z3T� �y��&�q����- �|����OV� 3A^�ȟnN0�6Nc4j��)��h��y��r6��}`u�5Jv@r��2��=#�����"�x}2�4{?�V>r�A9C*u����������~.@V�[���6B; pB���\�z�� ���+�7�̏�42�4�����wq�VHK����a���o����ü� �&g�Q�肾�^����U*�g�5��p�p;g��m�Q���>���nP�c?p�-K��^��+b�[���k����?�"���i�H�_x�DFG��~�E����v1�1ހu7�����=斿Q�eX0:��U�J��1 �f5�Y�d���b�ԤN�c����t�TuaS�q�ՌJ,��Pp�����b�1�ֱ���\t�x��t��J| M��n�q��C��J�T��)��[Y�?'��7��/I�&��F��*�?���<�򚛆۾�Z�e�W���V����0��*����L���F���Q� "T��"�7��_����K���8.Ĉ�������3�/�<:!L+�l�o�r�do:x�A�����0
nW,���4�����N(��ܖ"U�� ���rNua �Έ�@ �.�E��A�ͫ^y�V�mTg��iq% 7���<�I�J�\r���w@N�K�oR���U�����o���uo-4��à���-~�ߌAHr����_��º9�S�Q���#�����$�T;��Ț;�pZ�N!�<;_i4?_�g+Y%�������6�(��C���cv����������ld���GTƓ��.�ai�5/�o*�����r��O��V!�����Л�kp��s=C���^SR񥽠}�1-��J:����C(/�:=���Vy�W8��R�TwM��]�|�q	´���Q��5]�Ts0�f+o��>���~�ߴ[���B��D�GD�+���}q�	�a�G>�)��#� @̉�dEѶ0A�E�i[��]���n���U�s�em��&��]N0p��s�7�!j)<����WZ�6��d�?+1��������CaR~;����'�C�(��*ɳ�{�#$v���%�=���}���%�T���/l�i�}t�i*���Ҭ���4v��ϑ�8D	��g(��<Pi��4T\E��>��7���N�hk����g��TK�����FG�����6$��p��D����Y�������+��U��4~��(�슆C������2m��d�5�M�`d��x'�j�u�@jYҐC�-���U�9��6F�$5���u�nx����Y`��ԩ�޵���u�0��^;21@=8"O��qe��.���g>q�YEئ�2�
�u�NP���� �9q����VC��;T;a����G؇�Rؠw�㶦M|~���^ڼ:z*�ZQ�-�BW���8�:m⒁x�B�m�®�b��.0�<�~�ѕ;6W��yMrͶ��d���:pTj��r甐�Od��_4���7ݧ,�-�|ě����QQD���#h���c;�fW��yn��2Beد]�^+l#_����o2��%zJG��vQ|Gi.J�H�`E��k*��d�I�L��;"}�g��}�9�\M�Θ��0��d��Y�]9/7�Z
\ە+�;��)���\��GP*p�+D���4���d���Cх6t&����/�������R�?ѡ!�����&<ݵ/je���`�i�{���
�<�D�a�7��w��H��ۛ�����(��q5|#��z��o �9M�{^-̭j$b����a{	��e�+}=2����[3�����1o�Hj��I �9>��\9��|_s)0B��+!
Z\m��F�s�;�e��f:�id-��'��"�����E �-pH:�$9a�oK
��c����-�2	�"t)�z���Y��L�������x�|s�!w�����8����r����e�����(�̳�j }3K��[�{_�G��M��ו]�b����
q��k�o &�f�5�X�!��ߔ�>b�s�hK����ԗ��!��L@��/);�슗-�N���2���S����ҶP�+�6\�o;l1��f��������c`�=�_����?2��@�Y�&�S�S🷭eT��QdB�AH�W�U7�⡣䅔%�-z���#}9�2�����(f��������ek�7*s{����EQH��������z� ,��v�[е��;��,�eG��++_��p��*G�|J\���Q
a ��I4�)�p�G�)Z�E�u��/�%��Q�� �D!�
S�/#��ٔ�_0��7�0!c&CR�ʀ�3�7 ��(F��{ ��]rC���Oзj]�{�['%:`�ݛb
*1�ڍ��ܐE���kOr�c�܉x'�tF��d��He��`�D�Nȟ���bJ6�����􀈳ԡ� ɀ%�+xo؊����ƹA���Z��@���'ֈ��f6ΨQja�}m�1Qb*g�V^���j�d��y��yg���Q<|�P�
o�8�X���� ��V#��h�%�ӁK�h�Y^�9UX�/쥀�G�"�h��x�h.�� I��6��~��9��.2��T��������*�UU��q/S�ȽK�g�/��^<2P���C%�.��?�@�d?-B�L焒��1���Y%4�?:��܉��:p��+�D{�^��y���F�4O�c�5+�&qMZ��VO=���ʴ3|��"ᓀ���f_yX%�D5F��hYv�J�+�̣PazQi��fɸǺ{���H0�.���`&��z�-:cn��;��~��|��Z���+g�W}1�ʡ	��͐�ζ�PaUp�|�c�ȣ
�^�b�,i	�ĸ�㆙ڹ��q�X3�c3�Q�f?[�äi�y��	 ��!^=���l��b����^�3�%�i@F,�ǈ�?��(J�a�J������:o$9[��O)��O��*u�B�m���D4+��X�=��R�����̾.'��\2@�7�]��I?��-�c�{��J�]Ά�NM`%�9YJ�������?/���UwW\���/��Z0��-�M��6�?z�J|�g�A�1�Rj��m)��%������F<��ͼo]�dҞε	�L��,$�jy<~��׃��S�o��z��E�������Br��i��j�+ܕ�Nq��L�5z�rDP8�����i%��|NF����*C�e'�N,%�+QiCJ�]o1�di�T^ 	>���\�������\�-O�1����6C���o�R��(���j�B̭���L�g��"yCQU#�o�orx�U�N�������*�U
+P� �kK��R�%M/k�V!�K����q�rO�e�pm�2��|�4	6�yh;��
��9aʇ�F0;gLj������Ŧ�ؒm�w:'�527�����e�y��ǈ�c��z��n�t�\om(#Ȅ���D���q��>�,0�n���+8�Ѱ�t�U 6�R�?7�Y��y�pQb�*3���h�P�����G�B].h��ʘ^���\�ӻ���u����%Tt[#3����*iX��̀/>{��s�j|
�)��/Z���4�xk'�?����M�OV�F�8ͯf�ֶ�K�*���R�������-u��z�b��;m����Y�j��םi����b�.���)�B���U�ݰ7�ބ8�H_��p�Al�������-�>�ӥ� t�V�T���ҨvvL��6{�X�/��d�J��-�n��C�A�J��Nd�0���\y���j����<��
�V`W�q�4����+�'���"�fV����*7c�)E�bI{3o"��I!�ԅ\ 	�E,��ddIN���&o�ќ9�4�&�9�Z{lt��ij�MԸ��VN�����M9[���:OE�^�������U^{��:woA�AN���t������3��eq�&�ygZ�y�;����A����~�%ּ]���Y���
��1-���7B�9��@��5.��qw ��1#g�����	���OC4 �T�	{�v#�Q>J+\�*v"������?!QF�ާ>7Q��9M�r�\ 1��.Wj�z�p�ز��&YX"���q8DÐϸ`_����/�`�s�/�;�rX`�Ǉd�	�9#�\2wnԣjݽ�7';�x�N�����k2\ �7qhJ��=RK����F�6���t�d��5 k8�y�N4�޼�����f��͎�dd�����iUa��ӣ��>�ƥ�_���'�.=\�����(�<�>U���98/���-�ݩ<N ��<:��א|�*~�.����c�~u�YE�/9�}��h�O�V�Y�Wg�f�tV`�EU�{����7���X�yC����a/R\��w<~W�s!��V�m�q��QÐ^P�?ay�7�.,�Z��R;�l� �csʥxq��N g0�!L���IIN�L� ������3����:o<�ЀW]Y��O���� P��)n p`ɸ�iqt촏���.�Λu3"��\��zcek�����Ŗ$ҏLc;Z�Xgg$�v�ǃ�a�׭*�I��W"��+}�}����G�+=�-��2�	���蚽�X	F-�0����>\ )9H]�w�_��-�����JO��r��8P����k
�[OZLLLs�%�3��xEݹ���PH��as��pa� #���Nv���ՆT��*�Cj$Wy��k�@�f�q�"9XG�{�xc�b�|V�П2�"�=��A 3Ɯ��3['T���n �+�-��k��$��� ���wB�d��M=qZ��&��
���D����P/���0���םg�C��6C���)F^��]�T%[1�����b���	c}��p�E��pR�Y�:Mx<�7���O�T����:2>�@b��eJЯ}0��қ��
�'�)��8(�[�ǋ�4w�K�2�t�$�ǃ�.5e1d��Dӄ��E��JF����^M6"�5�Cn��(`�j��GH��Њ�v'A �m�6�4:��>���%�HN�-��]���ҡ�{zh���2���^!��͖1�r�	��x,d�����.=�V�U����u��K��}݀� X�t�HU���S1��2�U�`K3��:df�R/��*��8�w���qa2یI��1��\��o�Y*f���A�x���B�����C#.�7�s+����AW���ucU"h�oi��܁uU�����w&��`Գ�qզov�/��xЛ���g��,Yb���uoBT�Nį��7�{�����v��W}Ҷ"	,�jy�Ф:4�ط$4��ܒ�j�#�eUA�7�1͖M�u(/��|��X���6��N�-���xuռg��c��q;���en�/6�o��lz�ֻ��)2tnB8	8�|�?=�%���ƪ��Y,ۂ����Y���h��,�W
;Ɯ�s@p�X�4� �����F�.{l=�Z�w�"���G�=���E�R���L�0��n"ժer�ÿB7� �4��-�����!�塦��#�k:�^�/�ȟ�BOu�F�y0(�ČάQ�t��^n����g�a�5b�4/�c����p/R���J�^��2���yV--K!�_����z�:���Hr
Vy�Gٛu��0��瞊�z:�36��C�U~�C���B�8M~�d�ή����y�bi�P����e�xi�S���kbf�a��+ݨ��Q@�7�E�3���t�u��n-�l�q����mϟ�Y�qq�a�E8�����hQ��w��:��ρ����e'���|X`ɪH��ǩ|�)8-'�j)�=�&C��z[�W�@�� V�/�E��	aIg�(��7�M�D��A_�4��3��1���>�H�7�8�e���wM�z����w>ᡵ�=���(�����F�8�7ZY�����8ȩ��n��6?�����.��iL����H�Ƨ�H�����34 ��ðNM��S�B�bowB۱Ԥ�X6�D�|��=v[��TJ�\U��H#|D^���m��y�^��	5��٢_��_�c��[�"K��d�X�)��P"F��̷�z�3�^/^�Cy̏~�c���O�0���9'7?|ФM�d�S�΅��7σ��~���$�Z���2g�$����up��b���Yo����Y�BX���c��h�y� �ۼɘ�Y��Y����@ӊzL��_� ���:%�$��s��s�`����{Ī��;�B�0����B!��(�}��v�s�c�[�Y�o� M(�1HI:Q�o3�m1�����I?��jF�~���c��ٜ"��� �a,���U�*���|��2%��q�IP�4"'��+L�E�z�c��+\5�hNE�a��cr ��zG�ARb�/U��`N��^��h9�+QQ4(�5|�SĦx��Ry!9�}R^���ך$�uJ�S���`�-#�1�ѷ��.Z^i���P�-�
VG����6qh<�P9ȶ�}]���$�1h��=,�^aX� �����UiaíP]��Nz�7��P��\}P<���9/,�+?(��&�D	2���-��2�xN{��Us�dA��2��by4C�\;%OBѱ"J������G����?#x�|�=⶧�*ScgNe�Y�H����^���!'00����Q�4�F�U_�A0�Y=d|�l5s ��-�{�~'h�ò#��vh]���i�}i p��?������iFA3�g��ڄw+Q�8�"j�e��"��id�N�F"24�{�}#>Qd��+:S4<��c��*�Y�4�@����hvplT}�)7]�L]#�%�#���UA��Q�[�&�8��mz
G �;b�"��e���s�F��{{��/��9c�0�^E�;��,Ӌ�N=�y�������Fn��B`
�����J�"�3Hz����[��k~,,pR��SA��\[ <Q.9\���qŽ�N�X�O'}�4���3D�e���9e��N�����^�F
om�^���cк;i��>�tٸa��0��A�q�	�-��2�JXŗ��{�~� 4N��ߗ���wY�[j��rJ�Dt<y�B02i�2��n��7d��n����mv3!ˌEn	�}>�����j����ݒ-IG	
Y���$o ?11���Q��[1w�~<�$�_q���Ua���n�ğ��1��O5���V�!���Z�G��yp?m�1�8if��Yôu���lԵ�.��%��1�?�ʦ��F�V��A�P����ӕ-��7�ɥSY;>bd���k(gDoi����%s3wE2�5۝m��Ɛ[��:7wO k���5cp���ٚ�(����b��P������l�U�r����B�W>�P�K���E )3�# ��L
�AZ7>r�����Ԭ,̞Ņ�;}`�W��L���hLa!���Y�q>�XN��-!b}�@ͷ�yɱ!.��Ӵt�Y���e-nl9��1[����`u�ta��>�����R�7I>n�~<o��M��.qg'#C�xx5l�<@N�#��I}3��ԏ�9�;Gk�
C*���k��� v^�bKĕ]nn�.Ѡ��F��1Pg|6����NU���d��q�#�f$�7��,O�M6�޿���kQ����W��7L[0lY�����-YEm�B���
��jp���
���!֔R��ڋ��-�\���	�It�ཌྷ���Y]V���]J�%�GC�H��'B�M/19J���;�! �1�é$��5�P���Z׽��VGx���^ǽ�����b4s�tm�j��ǯx��0^Ycw�w'wY�6U�ڱ�6ŵ�)\?����X��Աm������9F�U�jn5��79e6":4�\'P'�ę)�88ޕ�C�{���i�4�qJ��g�Zq����$L<���-���e��O�s��^���O+�tX��0�p%�=��fU�a��FJ�t����2��iV��T.�o|�}/�:��S�s±�$���+����Ҳ�2x������8P�����}�
g��e>;��y��#���l�T��-�S���OAW�Xhϻp�+�
l$qksm�w���Q�C���-JZ���fs@@�����?�f�1i2O�M<ئ��o�,`�rОYu��[Qn�$��6�'��',ŧ�Վ.���Ԉ���f����6���x�7rla��6���	咏:���wp��Pkq�/�r<xd꓃��������[��y�:D����p�<�%�-���˲��H��D[��Щ��������|"����PO���
��e��j�R�2��M��f�Q�H��IP<��@��KY��F@`�&�mKi��lkf=�}Bϰ��7c&�V�&/5���jn�nB�O豵�3M�yʐ�t��N��v� &�-�"W-1��e��Pus���M��X��j��-�L4��Z����xnI�sz=?$u�8���89�����[B����.�A8诎�M�����݀�uU\$�Z$9�%���ZE��D�I,�lN������$hnEV$�2�������]z���!��u�&�lJ �6y�,��MgLz4�^�/��7Ҋ����b@JO��<5�/����\k��s�!��r�0���?�c>�ұ��h����q��}ԏk~�	ń��%��������XIm�׏m����	�Xƅi�`B=3wf�Z��E:�M��\	�����Y��-��h^�����V��o������:v��4%��F�W�Rf�V�����[���Pԩ�Y1��e5\L�f!9��t�Ň����5��|Ju;�A��cux�h�>��M��m"���L�v`U�E's��濿H��U��Τ�KO@N��£���M�Y.<� ��Q���}�{oS��6��~��jT����)�؂*9��r���F�ȴS��o�\;������ʴ�q���}�a��3��-~���/KZ�����`��(�$,��O{�8�Γ�W���} w\g:x��>K�����&���V=J رA_�����K5�Ѳ�_Va����ϱY�:��{�ӡC�^�KE��+N�8��Z��0�s�΂��������({����p�q
�W�@`V9k?���O��쫬Y��VG������ђ�aYZ�ǆ���rb�:���?�Fb�cPDQ���6�7����E�"�gv5��9ߑä��+04:����Q�p���;�G���2	�5bP"~<�w�Bsb
��I�h�֕Ύn$�#@�;�1�3;Ӛ�󫬡��^�c}����p�g�Xg�B[��N��P�0��ج��h��)[ڛq�3�Y�g�\,��V%=Q�.q��B�9�]=��挙�D�X��0�a
�q!*]U���o,VJ�8,�� ��K�l9�+���OY�NV���8@gT%9��M$݋;�#e'y{��}�Zc˾�ԩ�{���o��JB�Ή4䶾�#��*[�g���X�ࢂ�y��a�R�T��������.Bt�Cy����]����&�g�q�]ŧ\�2�M��Қ)�jg��HUP�Q�~β�y�H3��\�K��0I�;����e���E�d��i���ӆ�`3�Ne���8��s�F�t2?��h���KY�`���0���"ʮQG����I�P���Ii��Og�&���#n�@.�Z/_�<�3r�6�z���Uq	K�6�%4j�����ɏ�kohzWu/�[�~t��+Z/��q���+�O2:1���eb=��c�`��
aw"O�j'�݀�a�w*�c'?(�ncY���w�OmI��Um5�n�yf����Q�g`�H\xI�Ps�=Ğ0^ oAH�-f����o��YH��n�d���*���g(�w���ei>Η標��G�"���q�i?�;��~b�0Թ�%�����\4��G�MpL'<Y ܘ Lg����NǕ�o.�Q��Y�k��T���/�"{Q*; sx�7,�-�{�-�b|�3�f����he�6��_��j���<CL�c_��u$��`� no��U������¿<:w2a����tڤ��Ӻ��-��Nf�z��8�sA��f_���1&��@rK<;�?�4F�� >
�sԵӣq���6h7tE������y��R+� ߋzt{٢�rcB�g/�0!�ο��z'�M*TC�9�	j�1m��Q�5�\S�Ѡ�*^�X[��^�k L*�Go�����ڥ��ý���wRh��D���-*���_�E7/�dNw �W {�7��:�$0d�g�c���*uxC=�݇��ԢC�@S�H�!!̰gS�?Lش���Y�xg0r�#ۂ|wct�B�	׼��^��璬\ű�\�O��'���Pa�V��£��\u�|�I�	��5�L�Ce��~Gv�|K諭�7C\�v��W��0�ρ��n3	����Q��k�6��P{�
���,`����$	1a6�8�..�����~�~5mq���E������"�LB���x%�����@�̧u�g������� ��ˤ�g���A��y�T��;6�D��zP���)���T �=�������@�'���b���:-Q�lے�	�=��Aw�l�H�����Ȱ���hU�n�^��·���-USͶK�L�������#����k)���v.�P��^ /��?�Z���D�2$���R5S�q�{s��-�V�y�)�u��F4��q�d��0ݓ]z��5�k9�:�x��L�d�����<D�=����9��nφз½�͠'e����ĝ��+_mr�T���(!w���WAf�q�-G��n���_=��N+������ hڜ���Y��~�PGn�No�m	>.��q��[x�#�k��g�]%�6���jru'�w_�\P�v�h$.F�e���ọ�W
�S6F��g�L� ���'�[.�k��q�v3����&�^�R�+�'�j��иZqf�ސ��k<�+������}��n�p�㶘���F?�ǌ��9F�B�"��@�K�2�1�J�����c!��̝+ٖ� uB�7B�U˚vD��h��Ff�;��ԕ ��Y�����.Ney��C=�P�%e�R��rH����e��Vb�#������y��b�z�����4P�����M�@�C[�ÿ�	����+C���+c�%T��8ڛv_<�׸���}�P
���=pj٨�ر!���3y��Da����5�H1E)@�ƭ)2h��Ke
%�l�akщ{}?B�ഭ!R��.�
��*B)Lgn\������#�AM쐳c���d�iaG���r��T�ȃC�As)p�����S[��;���5"af����� ��(����LsH;�DU'�١�kS�U����������L�l�l�M��ϝ徱��?�y���X�h�������K�!΅�Q2n9����W��
�����B�E�[�p�6�t�^���y�e^U�����+��,�|5m��i�xP��t�+1.��@S�ɹ6�hir)Qj,k���P�3��F�ȥ�����1���$5��#V�Z]���L"m�2_�ojwTq׾r\��xrW�:���Ʉm�_(�um!�]ȏ�`��� ?=�éjZ�l/���?��� �QU��'s���K��9�}�^))�� �S�i���x8\�V2���d�����Ze�6�{ؼ��΍^=���Bg�K�V���z�k����X%��Џ����T�Bp�L<])H���+�u���ի��oRU8ʎ�EN��D�P�����Y�O"�2��d&A��
����e�����H�����O��,7��w�npO�D"�����Ke�9�d'��Ed#���8���-=]��{I�<Y��ÅA"Q�o�eMN���O�0M�a�6��=���ؓ�:��$8s��g�VFY�}5�͎������Z�Ɲ�t��5Ó�NÏ	�y�|�g~v��x�$r����BNLy��ˈ��dU���3̲(������}��Y�%L-J���F�a���Dm&�b�}�)�'�ú�$��ݝ@�m�a�ܱ�}<h���YW[M�"��]7t��B����4�e�X�A�t�}�t�����p�Tc��*|�ȉh�e����0hq��0�h�~CAur��؞��k��q����uWxk�*��TgL�d#��u��]����˒�9:�y��|�%,��i�O�#2夀�9����xe� &�g/d7M4c��H��{r�m$��	y�S�� K'��%�T�m{�?%�A` �-0&���ЕZiP�-��$:�x����g����}G�`��p\�vT�#�z�]�w�!�rGSB*cK�4��K�\�s~��@PH��bw]@'y�B�,�>����z4`�O�
�]\���@"���i�8����s�EeY��ĮX������Rɽxo�ݸf�^�-Ҕ<JrϘ��PN�MX~��\��,o�Rp0{P?�W%1o�׸��d�,V�/��\k:�7�D�|q��� 	�vvF�¾2�Y"C�{Sz�'b�a��x��?{���ʵP�e|&n�.��:�{�Z�Ph�!��i�����|9~�3�)�z#俱 ȫWM��T8��~	����JO��p�V�hKّ ����2/��>��A�|��/��Vz3�i`��S��E ���q��*[���><l`�����W|��a0�.=�	:��3��܁^fΚ�pѐl�&U��O��4����z�m9N	�ߺ�-��w�/��� W�b˥Pb�q(F�i������WY�=h*Əg;5v��uM�����9�M	܆�r7F^&���K�fb���{ ��K�VH{1
�7�]9��U;�ʗ"����h��kk��<K��#\)�;Ԇ@4��e ���s�k`��^W�d�)f�a.�;�ۼ�T�����e�o=�%M���
m=\hGBY&9�����Bcm�*U��x a�?E%�W�h&(��k���%=jN`�g9XV��~f�S�@�:NM8o�<>�՚z�epa����,���	������^�L"	v��⬚c���* X��{����_����A�2�yK~b>��^.牺-Đz����f�^ֶ͔���Y_	AUG��Y���-L*�[��������)Y#��1Ү�4���x����i� n�ۓ��I����viC��Df�S��y�uK��Q��:��k��v�ûƯŪ�:Q$�z�K��h~�8����t��P����l�`a�&�,�_RniF��o)GUQk'��S�W�MFA�j�L��>�1�2S���I�|������㿿�J�����S��ɢ�t8�� x1ϕo��u2<��2E�c�	@ٹ�uI/֗��w�!�1U�Wk���&n�CvdG��|��Y�P8��&�.<���mo_�� a��/h 73T%�*<؃��iL �?������m5�[s���M*���$mT�H�uΫP�!��;^���/����!����.w8�Q��TC�.ߑ	��o'/q�݄�U���r�m~"�v��6���D�N޻��$E��0[:�1ԉr��ߖ���La��f\Ù��0�ֶB����fS?e;������p���f��6��B.Gz��𢋐����\{��� Ғ��yMD:{L�mR�HapUH�3���v7���q��l����,6�� �6�1�W�[7�y��6�S\��ܦ����}	nf�n|!D`� M�ck��aNN�c��`�=��m$�8i�����K���(��=i����?D	�eHZJK��������D�=o<��<2c�������%�J�T�w�6tk{����]�i�m�7]�W�$ɱ������	�R�S��{����LZ�\�p���"�lms�A��EVl$��R[��"omȺ�1���=4�'�[U�A�ei�)C��ȴf���W���g���V�3�M���ŠRZB[�u�/�,��qo -��&��{4�*�XH�#gyo�3�����𚞗�oC!�i���7�+�4�%�s�Ɛ�Z�8�����5�[X$�L�N%�c���]�Q�K����פ9���P�x����/�����D{��X�GlS�~hRa�?�!-y⎛����MD
�L�І���05�'%���s���!_3`D�����.�%�b)�<rF��"J�9��#�z��$� ;>�P�bYҤ�R�'����Q�!�Hj���H��z�}}0v�\���/����fN�zV�=�&�tT
ׄ�ή� t|p4�z���v^e���ِuSM�����D�WH���%n��Dz�T7o�|$��bwT��[P�V<��Ի�!YS�A F�7�1=H��Y9������4�$��L�4��z�Tω	��w�Β�q�"�	�7)yJ�{eŗv֒=����j[��l_�86M� ��(��[7\�$s��:�e)�ZX�+5+�@r�֒7�	�M%F4�TM��ǚ�˃V|9m�����A�T�_��Z� �"� aG�(h~B���`P���a^�e9�/���D�r�������V���0��5�X��EDh�q���j���w��$�ɩJI���-����Q�i�)������[7tWl��n�jŏ�V��C���ၦx�r�:� :f��\���`.3lk	�����ae��7�X�n�������~�$���/����9*w�!�n����dw���m1͞J$�-�$U������\�c*nN.���U����}
5���]\�,���k:u#(�@]+[m}�� ~Ρ�"�&�l�W��i0�M���S�	h#�B��L���huZ����)�>Y�|iϪ�h���*Qg?�)�����/�OuC���*��"�I׏����/��׹��,��$���{���.�̴���3������q���
,����輰����]��bCɱ]s=��6�.��K�����l���bx��B��dD��v�d򡇒¿ T����X��.l��s���ˏ5��S&�m��ӝ�#�%[�U0�H�މkqODkd��뉺��IA�J���t�8�lȎ�Z��6B�2D��K!����
]k��)��VYᄏ�٬�.�y���Ui����?��3���ŧ}�*EA���{P-��E��y�M�;;�RLe$���r��*��iGP� �𶮄?v�˞p�י�ը��C	�vC�us��� )@O�=��Ii�����:z\�I4Z�d13A�c_�NȤ��wC$-���Z֬���Il�v�\\��`8�~�0�ֹ�R�JF�	'��� ��(8�Ǩx�8V�R��bnMT?��k��e����Ԫ�1�tf%�ԛ�f�Y'�v�i3	d+�z��m~�]O�134۠��JE��En���H�q�h���B�=h�W~����wK�� �X� R����T�R��90�?�-8]�q̜�Ħ�l}oǿ��*��ҥ�JR�u��w�/W��oa0�OZ�YB>ވ$�ﳸp<q��e��@��<�&#�ɥ��bs�/@�b��\��q��c��*a�Vr���F���_D������-��+���7��/8�qb��f[�V1J��oS9�_�
�[	:�}`��cY��+|Y4�^w�g����~��eڵKQ�r�@������GgzS����!����[Z���:�8I�Uw�5��r��uF&d�c��[�����(*���:�\�."�cN�vgV���:p�˹�7�A���&~�M-�*�EI[�[�<�3v��z�mm��l��q/�ÜE�Y�d։nE�-6�W�mm�RM�(����(0%�бgl�pCfid�d��]�� ��8 ��iu�z�҈z��K���9!I�g#�ȿ��9�@2�C#�e�r���pH���N�1S�+���yV�h��[K��q'n�]�#Je�a?���1�Ռ��>��(�ڰ�By�J��F�����)�o�	 N�x��E�MC�����l�x'p���[ǚ�^��V��Y���?T��� *�F��AY�򘙰�E�I�簩��Ո�covBǉ�[QN�Z��=e,�d��n�*n��e-S3ӟvj�.��c6oj����W&�&5�넞'���	�P���A�ձ��h�7��	��Uo��Y��F��	JK�{��n:9_�7�K��!���Yҧ^I���m`I���m���Ў-{q��c�j��D�
��ȸ�I؁�s|�͞D���<�?�e�T�V�Ѱ��H�Gvgu/҄�W�}x���0h}�
g�)X��d�S�TX~���`��� t���ͺ[���b+�F[ɛ[r/� �1��}x��"��R��V��U�����y��Y�U|�WѬSa���/Ei�����\-��
��F/�����OUB��N���r�To�A��rq6�cs=��Hp�HGY?�V.A��Ƈ� ���<��>��a�&���tN�H�� a#)�z�6�C׀��=$Of����p$s��<��VQR�w(����'?QW�����-��t���y":�^����� k�~���d�a�Z�]�ǝ����xI��b�l,�t���G:x3�2�ћ�|��^���N�P̸����T���\ܪ)���A�l�k�S�<�+G���,B#��+t1�%���	d��/ed��[`�曦�R0�#ua���ct��o��7@��ߟ��H6� �j
��/"ݽ�sm�Ѻ�qn�s􃼀*�̸_@Uޣm�1���#ė�><LIKUf�����0�No5@0�_~D�K~��҉y�dD������;�­-/�/:���
��	"�Y���u�B`D�D*�����p	�C�T:@]����oе��4����v����?��Df+��8M:�*d,t%�@ș	4�ͩL'4�^x��R�Xy�v��h��Xs��Z�P��}f���4k4A^�����o,�<!:����z�>�X�j�*N��p�iK��R[�q��Lr�S�2��d<�Y�c2b����o�|�G��|h:��Ag�#���'��"�^�xW�sB��5�a�Q1�W�ۑ>�h�?�{�o�RO���U�	�?qO�YUh.�����;&�����^j�^�s�%ӣ�4�-�3�\.T�`�.�E��2����)�G��U�p�cg����|�I�݆v�r����͙�-�)�R��N��F��V���R����}k�C�"��ɩ�p�2:�����7�D6��|2��1�^v􀖦�	��^�c�v�8�5b6]�)�U[�c�3������{U}�ǂ���(UM"g��PBIZ@꩛��ͅa�}�����͢��K&��)"'4ER�F�YW�.�%3��"kuz��E���.(�r-�*�����+��#��;�M�f�-�T��`�\EV�0w��c�"랃��E}ziR�\���G��U�T����� 6��hp�|:���kL�ȶy�W�`z��6O7��"�/�n������I+[v*M���`&H��2|�\�	g	���s2r�����wH�	ߖu^]����kD�r>���{v�?�)~_:7��=����_,��g&�d8!�x�Ź��s��%��b�{H�PJ�2�Bon��L{�!�xlƈ^���d��DBJ�ĉ�d����(�9C� ���R�r?���7:ϕ_u��������IG�]L��)b�����]�1���ʰ��z��/*PW,��a������
i7��ۇs]v�t?�׵ep�F���ܚ���U��@[8�:zɍ��c�x���P��x5�9��@9�o�W L��KS�|�3���;ʕ���
�Qj�8I���*�,�P�K��!�#B�`g��������˹��u/�r����2��S&q�	��� 絕&ǃ+9}ɀ�h,Z��F{�C���'F����G)��]�!�av:��C�ƚ}ҽ��օ?�!�j��8��H�x�b�Q�[H�IWa�3�M�S~πE"\�Ԁט����i�xzd����Z�W�j&�S�FJ1Nc�i|9��U;��u~��f�a���8�Q��d ¹�A|в�0�
Z�BƦ�E[/G |I'�o,�~'���U��a� ,�7L;���% �T��-�����f�ҴUCQm����k�N�I��N������&	TҗMa(XP�$�:��0��}�)1K`��H(��9P�e�&~�kLo@���W�}T�db� ���x@���D�;�ǁ)�Cۑ��Ҍ��5n����y<��:�Ax�7e7𔒪a.�$�$81����5ڠ�Z��vcx�T]�-(�[ԡ����@7�e(ʱ�p�+��!�tӯ�"ye� �����v��oG��ZA_�����=\5��y�O+_��{����(~�����)�-�`k�Q� ��>]Ӡ8������r��������}��6��"��`�y����8{P��\��\	>�/iVf�Q1ѩ#�>OX�5,�����b�� h��������L��J$�Kדc�`��eJ�n���y'b�2�@J\ޑ(�?n�����{+jZtܪ�c[��� ���������`�t���I�zd��(����C��ߴrM�X=������gis�	}lG�q��W-H[�g����!q� ��R�/������	���������^���լ��Jv��D^Y�'�ڛa��5�Hbߌ��<y��MڊOP�w��N���I 8D	#�����-a��*lFo��5�y�ׄ��|��G����"�l�5��E����/�ܒ�{��|��p-O�������c���쫹���%����u�)cO�f���=n�*DI������}�����;�_U�r[�A��<�*u��&�B���?�y�$�qC�^���K�+{�̢Il�n�>GC�@U:�J��7��F�^�%�����%؏���ض���x �Β/QL�>[p�f@�S��>��OD._��Q��n���1��L����}E��[�/q�8��zP�l+ǤGtʛ?��t�2ę�����
q(�#�g��Z ��|.��r��c�u�4����#��c��z�D����]�ɪ(������q���8�h�k���V%�A6V��psȩ O�Nc+q�� ��l���F��s��6-��lq�T'�c��a~����14a�呻�|6cǮ��֔���#��̌�r�U�=���L!�Y���c�E۶�
8���:]�8�"�-�dA�����i�����ϑ1���X.\�@K�t�����vKޢ�#��8�w3v���`|:�6��;�}я����DQ߶x�}��ӴE§�J'Hb������hIHI�z��5..��� �4x�e5����/�3���� �
{��2�%�g�߽�xC0�A6�9ع�a�\VȻ���θa�$Wq ,H�]�K�__��e.�6���4��� ��-
�i��^(�	OX�.�C�&�o\���:}E\�!��$i*r�x��/T���+��FyKH l)���ŭ�;�P����g��:%v[V�?��s�������"gI6k:�u��l=
ȅ5�2��d֬*ҲS��pH�}����[�1�kK����l�υ�{��$|�l���x�@�۴�z	�����z�Α������b�Q�rQ�=����?"�9�K��m�M�J�8��:�\}�2pT��p��w����[FÁÿ.�2C#/� }�NKCE�H�YgU��Ӈ2�絨��'�8������/�̀��<ޱH�隮/�p���4@9D��{XYy1��yq��l-���F?Q�9H�7T��o�D�[.�@����\�<�n<�sqA��C�l3�|�h����I`��BH�Y���4�g��y�]�+'���{Z�.���	��#�+�����Lq���H_����h�/r�0w��s�����G�Zyv�42��9�8�錯������Ž��������ѝ6`q�U'k%v�u��rsH[c�2����EEU՜�
�	2���ע �l4���mۆH�E%2�/�����{+� 9��<��r����:����#�ݛz� �%���\�Q.��툏K�{Ƣ�>OG�r�CA�YX3#2�M��j
$�"����@�%qJ����qt��Lg"��Ψ��_"����i�<!�$z�C�Z��R���%6�s6A�AԚƬ8lg( ��֞[d�k'��:�+�AU1�q��n-����ʈ�J��$|p� h���+x+���c�J��#��Z�3֟�zG�]�マ�G�j�|�Jt��vo�������]ђۉ��6�٦���$��c�Պ�Ƌ<��P)j�i�B�c�ݯg2�ϗ��1I�.�	���K]:�q��3�tf�΁I�		Ms\�:�o[��H�s9T  &�"`�[疞EK��)-���闒�L>
���V��K_�Z��=j���������9,'{#��w�o2�.R|�%�UX�9���E�1��Q��7�x��Z�;��6�_'K�`hb�������EN���ҀS]������50A�4m��	���VඕsE��27�!TS��EF�IE�v���w��Ļh�P�b#��+��C�`�5#��&�ѓ6���	�z�X,4h��hl�� Ɵ��UA �b��%՞��B(a�G��^��{�7�ߥ�/E�`�B��a[d�K�)zT��R.�H��I�8'��	�M���ǰ,I��m��Z
�r���Z_ﾠ	��#KYnQ,��|ǝ�N����L�-]��ϔ��z�BkU,hR���6�.I��%���0f��5�W�#�iZ��r%��Ja(2��#����RdA/�W,u���E3���]��-W��I�ׂk���9<���%ĳ�݌�|��-Bҷ�@�!T�m .��\�5�?�zk�*KX�ɤ�������)'��F�&߷�zM���Џ[w2h�'�&(�xt�*i��M��1q"�t���c����.����d�x�H*��:��J�v:��)X� ����>P��{��� ����|J/�y��n��Vs	?J���?������jk6*�!cI�7ɥG�4����"�y�u)ߖ�
5uB��d�P"���fR}��<�g�9?0��
΄̭'ɜ�U�{�F}�Ny�����#&�V���"gL��Wvt��a�ui��`���ΌD>��K6���|��j���݀���1�\�����o����	��n-d��P<2��V��A�~8���rGl�'�J0����p���@�C})��K�?�jұt߮L���n���}E'���S�@�p@4����;�bJƆ	kؽ��\����#�K�V>=<�;֑%�f�4ć9m}��j�S�G���/0�`	�:�@lM�Ҝ��5�247�3,��J�,h?G8p�NUr������x��ʑ�]��9b�A`��̴�7��ݳ@��Q&�3t�Chz���Ң�$�'��9�� �Y���z�m��u�������hW��M��[������t��]X�g��@�M�|��� ��eD�0YE�ȇ�M>���y7����O�'SN9��Sһ��lr}ݟ Pq��T�rbZ]�<�z'��|c(�r�Bf�!�� �.�1Q.|�U���Z�)�w'���֯�Q��A0){�&۝��eo�O4j��Jh�i�s �|���4�¶�Dx�qo��RU��Mg���W�-��zy;��cQ���,r�:���Nu�$iӃ�h"
���l��Ȅm��u����)UL���k-��T�d>���dh����
�K)I�x����zKU��CR �Q-9	Q�M������/�/�ȫ�t�^cE+8�+��z�s�rB4@�#�ׄj��t8�j9K���S>`��|�YP�,D�1ˍ�n�[���C`in`�����"M�-�/kV����佲&WXk)�q��Aȉ����4k�^s"��R�Q�ux�o��9����~�������]���4��y2eda��V1a{5=vÒ)#�;٧l&�%P{���f�X�I׫����5ɴ��erM �骃�Z2SaK��^�:�\stq���c�&�Qu��l*&%?�X�� +�zҸ�4�pg��g�F8����E��"�i�uM��(�H�ܤN) �K�'����~�������E����C*K��\L5���7��}��\;G> �M���4Uj���f�}+���qhQ�tYJ��3c��o�����-V\::�Y�&���+H�r�]�{:�\O��Gv}CSh	�������$$9FH�]�|oA�r��a.I�����	ʌ�P��y�so����X` ~��#C�+�̭=�����N����%xݭ'�>�+jÝ�pE��3���ou-�$�(���ݮԞ��w��(.�x��s�#4����R��aiƍ$`�_d�y��|>{n�{AKѧ��Q��6�t�`ʈ������F᡻����5��!�G�X�ɯ�٫�8,N>!�[ZPNN�dSX�v�4�;:$w�5?���&ש.h�� ���(W"@)����5���C�f���YZ�JSK�Sk���� ���m���y����*��м�4'��}���ع�A����+����K�z��j�{����WZ�:j��^˨������B������T�^�)�1Lw�}���0T�j���!7	җ]�j�Eҕ����?!(d��6�޼w�̍��Ob,.G���%�,ʠ��Y�7ޝ���#������� o�B/(ϣ����5�"ZY�
��-�����i�?>��K���c����R�՗�̙�Ed��`]�n#[Z!�2�Ru�鉶X�qqĮ`��&G�@M�8� ��(���gq`��J(k�6	�m����7S%u�8�`l��ɴ��D���R�o-9[m��^@{|	4+S�T�x���V��	�|~�Y��'��LD]+)��n�=�"�a�s���>T7�~��"viz�(�Jz���o����8o�QN�)9����:�y�Q�l�al��MOnA\x�1"�&�7��]���'�uj*���}'���x�$��T�h�I#W�G��2󳱃����c����d��Y�YYa�!�'+/b�Ԙ]���F�S�7��[?����>+FT��򲪤�����'�z�k�g\�)�>6��x%>��p cFuc����������U
�v8W�zK��l�7\o"R���FW�/t����L ��U�2a>���j�M`8��[TK�B@)�D�v�=G�m8�\$�Y�q��\�u�͎�U?~�.|%�T���`�qȎ�,�8��@{[1aLccKJ�C���n���vB�.�>z��H!-�A�k��O��:�ۓo�AoN�ٝ��IV�e�{O��i�3x�Z���#�;��O�ŷ"��XgxH���:c#�?7|�Q��B�J�q�>e��z�t������ű�<�z	�N7�h
ls�l!c_t�Lexd�a31���_�3�B���2����+8h�]/.	D� �X�k|���!������NXa �(���71I��a�w�2"����'~\�?�⡣���
w2V�n�9I�[� T���,�꾾�()����̏wY�JA�z�*��9~�W'k|\�o����~�/>�F�sV�l0UOg�iF���&:B�.~m:S*��̅�9c����t��'�Dk��<b�;��G���B�َ���. ��=M54Thtd�${�Q��2e` �3zP�*F��l����=\7�\�����#a3@*�t�f'��!��.�} Յ��=m�~)��N0S8_�C�������T3�j�V&p+�A�'�`�i�"G�w��09_����0��Z�j�˄	�ρԥT��k
�����r��j-�����>�ݷ]�8�9
�;}�/�B�O����@��b�h6���i�L�im}�Ǳ;X�]��&N��ȑ��+0���l��bf8�&��+��y����'���p�Y�;���.G���ݛ�x��ŵf�uN��	܇L��Y� �֧S0݇�ȼx����1k�$�cb1 �������&Q_�#��R�����y�\3�c��O�p6x2��F~�������깎���[i�j�<L�ۊ���?b�����q?'N���d��@�6�w`�/Ӿ����:����rI�º�U'YB�s	W�b4��p���Aû	o��c�UE��L�Y���8�*ti��ۻJ`�e��@��z9F���"�w�^<Ia�BU�	ֹ%��,��{��܀����Ɇ_vt�s�WT-�F����K$�����Fƺ��̵J���g���#Z���-�&����s-�
�.@�M���|�n>P�騂:E?�{��I;�HxO����~o7����=ك���	���)q��'{�& e>i�b[]��@����rgc糖��`��}�[jz[���
���h��a�N����8�u��IB�v8�B٪�����p����L�T��q4�EQ�t�G�y���x�Q7E!: ���j+�;=y��^0�e-�C�h�&i^��Mƶ�%�=�]�m�\�~�)��-�J�.��G�Qx�;)�b��fÝ�����<�p�#�(�%��V��5|@E�/gr_�dK��I_ևS��n��r��RX�5���kL�����������_����mI�$�wٽ�^{�ySL�)��g}"�`���{�г�s@�����)�CedFZ�kG��P��$�h�=��n�w.MwڌŽ����!f|F�8�of���\�ø��������n��_���ޑ��]_�~-I`�}%��{�ZF�c��3Rh4�z����˓]���0�A���>��7��b�e�B5�!Z ���ص�(`��κx�q�H'�ũ'�6���Wv��RB,A�����bL�ozW�͂�>(�t��Cc��e�@�7"\d���6I��ߙ^�\�(�����i{�k�dYH��	Q=��x�����?�L^�QYuD�_��@��c��B/���L���}��X�h�U
zF�K�ǻ�\5�tr����8�xҐ�Ǟ&����:�!�A��� 
�|��}0:�������Yޑi����Y�%���T>��ն�����s�2�| ��k�������//=�mT�ize5�Ӯ��5TĲ��ܑ�|7�9��ц��bF���Ds����M����
�|������l�>�p����sj��vrZR��xw�}�EF��"s��O�7�S�4o5��ݰ�Wcz��8L����Ĳ�VUJv2�zؒ;ƽ�����Ń>�"�7�g�72#8E�zr��-�bg�+�T"$g��9Z��	o=��[0T��� �19���륟�W@}b}�=��R��Q��h9�^T�,�ֶ���-#2u�o�\I�>GvB�q.ލ^�+`����4�������5�H$�k��ĤL��+=��`�p�-,9v_�;��m�)E%!]�?�{����{�s$D_e�蕻@�r@�]�5Eٛ�����v�ևX0W݂
聣,q�J;��*a�� Z��d����lq��wPS����D��F���3�=@���ul2�qeՄf��4W��B��A-/�ܞȂ;9��yv-,��?A\�0C�m��H�s�M�/|������&��:%'��z���j	$ �C���µ��R��B��Y�M��	j��o�́�B]���Ʀ���V�pᨯ��'�R�ƻ��.4)@1��Z��s�a}7�G�A�����7�j*;����QXy�֧�Y�/y�㜭1^�3z)+��*乫d��\�	f��k����0���8��*�uߠ�f�RH`^$�XwK6+��mM?03��#��u5�^�$U�|ւ$k�_�ά��������*��4O�����o�s����a(�U�KZ�8�4�C�ƋaئR��Yn�����!���m��Fi5�72���.���E�Nu���p��{a�p<_� �a����� ��QWǎ���S�(�/�g{Z�(�m��8Ժ�+2e�4���t����M�J�P��l2kMG�쵎��X�{KY/�:eH�� �t��o�Kb���Ӹ�␏� hᄙ�}�.�v�u[v�S�޲:�г�V#9v#{�,R� [̄�u��.Ĺ۬�%�A�V�}�&��9F��F���'�t,��5�Cg	�	�ǋN�~�i��܀���4�p�^���@j.��[��8=�D��� �ceQ�	1Y�噴�Fg���}��'�M�t���L�7w�[�g�I������A�:�CV�Rz�B��1u�oڲ��3��:&u܈$'Y�A���;���斬�!�)¼l�4\��_?=&�=�$D�b9n�m\N�/Ƚ+ō?~�^.@k43#Aw^v�rU�H�
�G�H����t�6��\��jimq� ���IBEb',oQ�u�z��sss�c_w����b�c�Z��a�����!�a�󪸓�;�r�E�6\0��skǵ���8�U�p����&��嗘���9�;q7��}�����b'��0,@�cĄ��*�<m*oX>ub�����j�O �궉�ݢC6��5^Jp��x���Ba�c�e��L�~���\�؉� �@`�ZL�`�}�	��ߧ�)�B
d�:�Y��R���׆�×�4i�`�Q��z`��tg~�ݘ�b۠޸�6�����|�p��Aw��R��Z�ǟ�%�9���!�Ϸg1�s(,�pn����Y-%��N�c�Cn�0�N��֕3X�e�: