��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*���� �]�܊���̚�T��]>K��m�\��}�"���uB�;ht��@���itW�c��p}v[䈐��!'�2L㧴���1ۖ��d_��e����,�}G� �:�xt �m%%?/ ������y�����8{7��Ų�2]�O��R�y׻��Rd���r�8���6�0q"����t[�{���W�a��g�^��dk��� �W�j�_R�i�l>gp��UG�Bg�Mk�{!����+�z��0Ҩ�^-oka%�bOH�ObP�����0��Q�@�����[R��;�������3��[�$N�c��r7�M�>pP��I��@hV����
h�8��l�]B��X>Y�C��LcΌ����""f74�R����t�<[]ܵ[ջ`���h��nO$��Co����Gm�N�!��/.�g�"���]g�|Qg+繭~�#��G<F�%/,<4��T���[�\�1%���S�4��X�r�/2�]7��'���D�YN��&��<KW�q�.�c^�I����2�l���(};����#���y�P�b�g��Bz�*,�L�0�P��@ $�]!�� /���c�d��/9�P�����K�Q�?�O'j�v�; �&I�n�p�+��6�����L�ʄiQ�rm��pY�ss<һ�a�%�4<�4��o�u�M��;^��gęT���cfD��!���V�;2�$���rc����B�v~�C����T�����Q?c��kjI�	��c�x8��:�{0�&S��x�tm�0 �t���?���%��k��[�Bt����܆��x�SN�������^.vC�IEmZ���k��D�����-�@:���
���:��<k4���� ����mW�Ωa��/�R? hQl'�?�u:p�30�'�'"�F�?�	�F o��,2���),�oU��!${k� 3Q�X�1�"[��z�k�nA6o�`գ�������UG\������ �A8����ՅK�EZ)��(�<%�Gާa�'����u��.h��B��=��دu�I"<��^7��M��l*��F�1z� !�\m$�m��ZrϭPN�x��P=2`��O]ś�m��\��M��p>*�uݭ�R�	���B%ʽmLͫz�#�NX9[�4��#�(�`l'�!>�� ���p�]���RO�qh]-f�i7�(���`����n�"�i�8Ui�L����i��.m�&2� ����i�{����iy |j�P�$��	zG�*"�)m�R�m����7-+���"P��#]a�B���;J�.�S;�Z!��b8(���H�g��2j��!��.W"�g��,v��]ķ���=��a�����u^��vf�pG��9�P�SW3:����n�	lU��[��?�>RF�ǫ��
r�t�VE�ڎ<��aH����##��{�&O	Bql����W��G���<��C�,k��5q1���X�1���Y�z.��=�_~֊�c]v�)��cQ��W;�t�ӝ���D`uvSt��������PKF.��H@;���
wn���c�U��6��n֌�B�O�W?B�|e��E?�x���d�R���ئQ���و�����in1���Cj:W�G�	׷O�U�9�^��� {/Ri�C}cv�=��9=��a$�]p����Y�� f�3X���aܛ�K��Y~7>�N���Րo`sB��8f��i����w��:i���W�cQPU&���z��Ւ�T3mj��e�ц�q��L���y�U��2�b�׮9��[ݥ9���/�� ���"�L-.�o(ǢI�8a2m������T@�joS�`�K�J������ig��9���k�ͣ/@��J���Ǚ8-�xf��?�(@Պ�TW_:�G^0�)F��L��眯���kIw���< Q1��R�߻D�.Ϲ��5�Ͽ2Q�굊�$[�J�ʪ�ƙ�?	��,��ܙ��=�}Yq��"��el	�"����r��}N����O�
�&��f΁�ʍ=�8�B�ɛ�.�a G.爗`"�Aγu�O�]�#�ĜMB�;��.o��|'�$r�~h5�#��6�kVJ���/���#��;�
�M���XH�+a��T#���������cmK{Q$���[�/�a�"�h]Y�4��|	r���c�"�ɤ���@˃����m���X �9�����')����_�T#IjbxQ���h�������n�"J�Y|�%��
>"�����v��g��LHz"+�GVFL�_c ��r(��nE���f/�\��Zs����MH�K���f�xɑU�J����*����x������� ��s͎�%��▋��k��K�)ݖ�k6�O=_���J�>M��W�_�Ylq�&0K~VD�Z1����$ťFF�̨�E��?a[xĬ��cc�N��_���v1�q�1�E�%�,{ iܾ�ϡ�oX�#O�}�ܭ9��ւV���W�W���U\���h���:9K�H��6���~�K�<'3a��K)�mY�����MW��������΁N����!H�B�c��/�o)4`�iՓ(�?�����LNM
�{��q��*��Y����}������F9�J�G9f㥢������Y�bf��.��&�Z��#A�K���x�UI����Q^��Q��pϩcexvTb=	Ч��B�?�2� ��b��c嘪>�a�tc�uԹ.��J�c$#*��A��,�Z$k)�fRCN}�d�ȷ{���J�l9P�L&�`���r�cG��x����**����N��ZO����J0���~�=�Ұ&W곳�#�ܡ�d2�'��z�PUk\�0�x���Q���W�m|)Н͠p��'ʊm�^�oݛ+~����R��b���r/�ف�Wx�1�i�c��鬁rr�p1��}nk<�@9Z����1K��B�8y�=�v��r�e`�z�-�L�}Z#4�nK�7՗����N�}���P��ȵEդ�j�mL+��� Xq��8;�xAf�>	�m:?���O4J~M�!c!_yGx0��]�^VO�/_�SO�I/9�AT|�=���kk�'�����"��wi��V�hP�>]�s)!�8�*/�m��_��3�r��Y""~�U�S��!���]�|J��@}޿;��_�\h�S��w��F&U��>���|v�U[�x:k&�$��i����查�+�!�!����6M�y��'i�Z�x���fŹ>����B�E����ҙ*��S�Fk��W�Ӂ	
�9�O(D��"�);�	�����=,�s��pm\��/�񡲸��(!㩀��T�r���¾��w�����K~A;U�t;aN툶��%o>C[Ƞ�8�����ܸ3��pq�������]�<q�EE�������g	�P��"�{�$�c��q�T 0�:��۬���X�����%I�!>@k�l?b:ڛ� ��B^��_&1ӟ��:y�?,�:v��9��|8/�72��";Е=�a��K�i���}b��34��+�l_0'��;۾TԦ �}���7W��BOl:i!u�"O�i3�ta$tϻ���Mʵ�)����.	�}�'�B�S1�0�eT~1 �����y�T��W~{~H�Ε�_��:<f?z�� �w�^>Ph�ӭ����M?9�����U��!��Z2��l�|H��Tڞ�|68)/{:�'���zfχ]E,;�V ���p�?טa0��m��oO��G"t谣��Y����h�c���RY2���O��` >[Lr�J�)�M�����%$��'�U'-�02��뭚n�\�2�G��d<cr�o�%i�*�I$0��E#6�q�0�R%G� w�wq��y!Qϔ-��-�Y`����K��`��#�@&]�(�.��5hۮu��̀��r��p~>~�.?��z��1�״������f�������"������C�	�h����`B�8"��Fwnz��� �C�v|��X_W��<�Ң9��Ҹ"�;skQC�qX"�N?��VA��(F$���5�w��ξ$t}�� P�S��J�8��k(��ON8����~`S<�l)�^-d22�͊��۫O���T8�Vk���$~[Nϲ���u��ӏ-��6Ŭ��Tt�J Rp&�\���H���PvF�mH�ƛJ��-i����B���#�l`�2$����
�g@�[�@:r-(.b~�����I�dZ=��K@A_-�a3$c�֑K�����s��1�Չ�l��fB��M�~Gp����x��r�B��J��&���z?�%9?˦�O�(��y576���+�4A�Ӱ�Z��_�Zq0����#���ZG�Iiͱ�N0�J�'(�������+	�u����Fa���)�Ÿ��0-@��|���}�ϙ;�6ҽ����*�@P�-�"L��x��P0c���y�>g�f��}H�
6��[����ۘ�Q��k���6�բ^7e�,�6)G��R3���fRͬ5W����+{��X�ѕ�O5�6a�M�G�M!��rwZ?I���: '�RIq�!�TgpͣR"�;c�����=��{��5��O�� u����8�A2O���(�x멎̜N���'8f��B�R�L��;�w�f&7���F��X�#x?@�7�[El`��-0���7B-jBveռ�JI/�Mt�GŭT�`�iT-fXd�ͱ+I{K�ن�~mu4�.�v�V���I:>�Wо��i�}�����ߖv�0z��6�}"��Cϫ�j�O'Qv�Z�i�5H�<��-�qC��p��	|h�0���=;EDT�^��@���~)ƫm�6��ƟWS��"7���vS�Kd�cb��_���lC�<O����/��!�!O�(�]sؑqi��\�[�6Kβ.S��E�&�PP�_�&��vDx�y�g��8���՜��ƥ���p��'=��P�x��2g���2���+������>F�N��b�f�(�����m��_��0/�;Y��t�4�`F�C�^.�	t,��,�d��i� ?I�.��MTf��h�&H+��h����`����k0A,!�������*=J����G7���]��ÀU$ I��b�Q�vQ&נ�/{5���-���˥�D�M��|!�ı���h�I)/�	��9u��r_z�0G`��Z�Ww�#�"r���Q.���P�2�`��'�Y���Mr~����ځ���nGP���$�g��͝ �Tr�������1
ȕ������F1"_�\U�#����),\��>I8��c�J~	)�����6�iǷ��(o���^���>�7g��\���ݼ0�.��EKBħ���z�(��$�bT�_��$��Q���CVL3�=�;�Q�vu���D�Z�
�yQ5�+#:����E�S�Y-c�����w�&zP��qGu����~ի��1TS�k#p��EA">�L8���q�` �/aҌ�Y.b|N�ƿ�ɧ�]�z��0��X��o���o��%���ݩgc2�	(BDx���./���U�
Uf��!ƠP����Ĭ�s5k8|q��Z���2!0�洿�/�l4;�MZ}��떶�6r�L��֩p�d<s�.Э,�C����3[2�L��ŵ�/���j�R�y���S��*Z�xy�;��j�.E�C�p
�����Dx,C�<R�������a��<T!�d��7�r�m�3N8�+���-�n-�+T�@�1�M~fgs;��X<L�`ha�!C���1�ś��n �=)�4�cd��z1�鮛��
����#\0�o�
4��p���6�Q�ǀ��J��1(W��}��2IM�i��SQ>Ԫ_�T2���z��#Y,
�Zx��	c���_�p,��v4����LĘ�����j���Rb~���e�"�TH�R��V���c����yw� ļ��Ջ?�4�XJ1��I`��������ʇwTů2fD��������[�g@ ��#�M)�^-!j�y	t�O�-N��hl����|�b�k�Ab���_��Z��յ�����5#'3��a��.sEa��3���Z�Z�NkyG
J\~���|��g��|�8����iT��X)��O�ո�51&"_;e|t���!�_��ʒ�h[�*�t��[��pJ���q'�U�6l��1�N���B���@imƥ�U�,���2%�ƈ�6Lr�B��PN~b>)�Gf��^�H��;,{n�$���T���B�$o���I ��Ť�F"�t�h<�;��sJ������֪��ӫTbX����p?���MS���ڲ�Y�{��	���SW��d�
�,�Q;��M-���a��rFDy�(���*�[��Z�;=I�H��N��䍀
dnjt�V'���e��
dH�p�>�p~/�ј�+�D֡��/T}�M`���#�h_6�@����`�`z �G�{�K�]=��Z�Vă���`֯be(q�IKZX�J�M�IH���7E0Ջ,��"�qXlm$$� -v��/�OQu�ͳ�W�`7�c���1B�o��˳ѽ�3�c;����ʢ�✉�n�kӵ6��A��h�s�}*F��c��g�z�v�����he(=����*��
f�L���_��ɶl����c�P���qދ����tm��!���CA�h)�@�濊50�&�D��K!ɴ��V�n��L@!٭# p0�ʲC�H�-��|�%����OTȧRL���Iٛ��B�C�U�&>ǥ�8���Tp�-L�s�W�\��{g�vb��,ZJ�qU�v(4��ַgK�_�m�S]rK�/�`����8����}f\����� ��#���V�͆ʢ��N����JƤ��0Ō����q��&d�F��$Vz��Gfc幦$8B�ׅ҆��8_����w�r	���K=wqR�����5Z�tiM#�d^͟Wd���lT��2bp���?MuL	Ý.�8�]1��<�������XF7�������B����S:��%w�����}�߇�iXָ��q{���/����M��ϓ	�����0�gQp�G�w�S,�H�G�m�ˎ�w-�z�y�ۙ�!�䐂�m�#��2����d����}��':��A:=��+�_� �n��hV#�%ݚ�.E�̩#T�&��/]m-�٪��\m-+�����{Qg����i�������_A:���7~�JJ����Hi����t����F��6i���r���N�}� �F�\��)O���HyN#�ֈ�����s
Y������"@�ʆں 4�'p��0d#�Dy��O}>c����)�ߦG�B�J�?a���%�Qе H� ��g�R��ǯ>��Lz�A] "0L]CՑl_��G���ߜ0n�ܼB��o��$�`������G=�Fz���5���6;=:��°���d����et$;P^�����8XI���D���50��%q�����2�\+�]�< �M�ʲ�c�J1*�}'9���w�ɦ��j�/C#����Ä�{��{yw-3r����%�a�ѓ�K���ı-�y�ܧ�Za��[���,��C"����Q,�ң�`���Vt:Q�:v����!9مT�IV�䃻�
8��op&h�}�/~���_�e�w��C�U����۾GK�Upk��^��pko��R|ڲὕ���-��?�Q����*����-�ԳX��c����j��k�-��e��n�4�2>�p��Ͱ��1Ӭ��S��8��P@������U��?��Z��������H���`�(e?�,f�_�Ks��W��lg �{��kө�5{�<O��xfq�^�*O�����i��&V��wP=��x����$A�)z�����,�<�)�0XN���bXO����H&	��V��"�������VZ*�L�jaZl%��>�
C'���+�0wv��I5�ڷ�ͺ}H�&k|쩽6��W��	f^iA�'ż�5�q�dZ{�:>�� 1'�5F[R����>���o�F�Y.JY/N�d�* IQ	oN��`�>� ��aeE�.��:I�{��ei�̠:�`�`�K�N+��h��][ٓ�8ѐ��m�\�������U���XPDp��s�֪@��E�z������Ԥ�S��uQ��$�-ZK�⤼f�j��r�]�>�X��J���^UU3T��{�T��z���Z�h�I����n�
�C�O!ӧSq[Z�����%���Qe�]R����MU�NĎ�$�i�Z�sX��0���$�i�	��e��(D��q3[醚����	��d�Tcz����VHoo��8`P��b���;���]WWt���W%��i3<8�X�x��(Q��tQ��TPE<N&ۛ����W��q6�\�@�3�H�^���ۿv�B�W�́��~r�Hג��}dP1��^�XE�V��3h������0}C�$sMG������)I�AV�[~�3f7�����_}@�Kq
޹��O�uU�fR���
�.<\P&0�L�[����;��뱊M]o-S2e'��
.�Mg"��B֐,��' q�SO�C��S^ݳ��K�{ܙ�BӍ�3��64ޢƀ\����D�ߖ��k\;'�VC�b���V h��..���do�b��!�$!-n�L�V�1��9�,��O{�?4�Ou��ǵP�y���4�4Ɏ `6�Sp�ծ�ޯQ-�\J�<�Pc��4�F�3In]��螜�*��[��^�|��)$t?�f@lNX�Q,o?�z`"���w��>����2S��Qa.�1��&3$���~U�Q��cg�h��rL�o�x���eD��E� �e������()2�(������{��åS�~m�n��0���#-~ǋ�5/GF|�ͥ"�@�#�Tec2����Tb���:���ڽ]�S�X!�hW/���y+��H)���Ɏ��8�R�<��S�V��S2XZ~]|��y%�|�J��`��>QH������z"c�E�xcpA M~���W�%�*�Md`{C���G�c#k)�߂���?��M�HGZV`�I�;bDj����FD��,\���!�=�c�����'?�ފ��S�2e��<��N� ̕3��Ɲ�[Z�'�>��Ñ��l�G�lk%^ԡ_���,��xQ�ϙ�d�i5E�{?�$<}�I�č|��v��ͯ���*�Y�iIm�Fz�Pc��n���G*������P���ń�
��t�� I�t=�����c��dn��0��Q�%�E����dӨفcʲ��8�(�3��0�gV\�r��yhT��Z!��M���A-'��k89"#&cO��W:?,�����x�� '=3�{�J�b�R�#�* �?��6Þfw��<�|��N��^2���͍��rԭ�^�o)>�/e�g)��s<��}��1!��m��5�Ń���?����2�Ǎ*�y́�j&��z�}ߵx�>z��1k_ k��#g�3���1���JDر���	���]��Zj�fT���$�1�k�g�R}�9CB*"��ӈCl�u�j��.h��_��N�b����W�װUtx��WbI����Q�(��9�>� �o"�9���v61�E����ar�>I]�V^�����A�O}��2�@�6�󛞣�%s"����6�QW
��8*wޠ�T�7�*`�nw�j^!�7��?��v��E+ ����)���"|���U ����)�s�I0�Id׏+�~l�cs��ʦ��m�TZG7��@XΤ��[�d����O���0�.a�loY蠙'
lZX6��}��Q%�7{K΀ �5_!|ٵ$Q������㷊}d�"%cG }������yo:i�����USὤ��'�s�{��l�>?���m̋��/,����1�h�:B�$z[���(&���㣣4j�2��`p>Ud�Pp*�t�@�� f�2�!������b�J�Ž�؜��*u���uz&�j�to6��(�m&��:XS��Z�򛂬�RRH+��O`�̅ut���c�[��G��ʹ��S���ܝ����W�
�B�T�U'.��'��c8��j��g����
y�s��<�������ؘ��� �ׂ�2�29�{(C���1�zR	�,�z�{	�� �0�o-��z���*�,��_Ћ܆9�`�+��6`TՍ��g�L.�⟟ٕ�������~!�%20�2O���x-����R#�T�;M��q}3�VW� �Ҏ�b�8����l�jw0
�qk�-!�[���k0g8^�ZVn
bv��\�&�~��H������V����f;)�l�U�85q�'�<d��Xf1�/�/΍��]���0�C� �����g�@�1C� �ƛ�ISq�+�NO$�Fb�Ϝ����)�5LqH�.T-i��q��-:;\�#Z�;.>�^ ����U�������Q�hYYm�`<�;��؝w��?ky$��_Y��hL�0�"Da�:焅�%�}�&q�����6�x���BG)���6��ۄG�ZԚg������̡Л����M=�#�����gD
�����:ΝKX�����6� �� []��4��
�#������y���>Sp������O���-�����P谯�G�kng�v�O���%�����,c��}Y�[xH�5����>�I`MD]i��s�٭ =r��|��`�u�5�ۂH��]KVg#�/�����t9��ɨ�5�>]��ⱙ�)����]�G�(������l!�/�`:Ɖ[w�Y*�%�mt]���U�c��)��-���kܰ��2���	!p1�J1*���FR%	ب�z�GuiM��g�M�I��B�`y? ����E��z~g�FRF�k����1�^�-Lv#�ĳ�g�? X@.�<񶾐���Q
*s+'�?��1�	ArH�[�oa�$~E ����!�h�S1�C{�|���(��
K�\�{;[�U���<!Y���1fx��?.ZL�r�i�^&YKs�����;e�:��LΘH!%��2cj�%��8�ԭ��	F�{|��Ls><�Z����]yԨ�.���!��Pʝӌ#��i����o jŕ�[�rS�?�-�m½��ADq!c�.��x%<Y��c�h�(/V�?v5U�3V�l���"d�ťVk���q���($8�j�����!\B��R��a��<	L�Y�I��ҁ-��~&EE�
���;���g�����*`�~&X\����J/W��ǈw�]JW�tr�Ӗ�'J�ԇ�C�;�	p��L����Ǯ�H�P�c_Ƣ��i|�_��i=�&�-[���D�z���uM�������� :h�ǫҡ�mIL]�X�\7O߫p�cԄ2�q��H���D9l1��27��oQ��
N�d�&F��{�Z�N1�IAp0F�i��g�oK&t��e�S ����lw 3%�j82j�NΖ��S���|��Y�xf,)$����/k�� �ķ�/�a��[�����}=%�H��+�<I1�"�f����	0lA(큀�j�^��u�pQ�����a�"��koD��xm��T�o�'VU�?#U�Ꚓ0�*����1e�R�s@?���^���j8�^�֓�|�B������2,w�2�+��%#G{A������4�� �!�+�lx���1w;-Y�)+���7iY��H�W���Y��@ 3�kM<��8{��wB����p��Z��.��=4� |h�Ǘ`�:p�b��Z1G�f_"~��A�L�����J���������"���r�յ01^�E�=U�eXq4F<�@�쾡U������,�u����$ˁO��u��v&�jC��x;_e�)v�f����.1�L����b�dV�E����x|:�j8N���.
n�"I��\��f�@����G����a�$hh_ʠђMuq�p&f�R\0�W����Cba�W%����$."��u����0���֝�)2���F�D�� �շ6T����?I���a�����3�2 Z��c�]�}��H\��6������GOy8H ����W���,Y	�u����N�,\ƌ�"�%���G5UѰ3�7�l��{fxi�m7�[��s?�	�W�!���<��v��$�������9��;�F�����sI�_�dS�ĠfiZ3O��E:H{���2�JI�a��!f�^�Ѫ��7�v}9�nA�$��)�)\��0V�"-�Mۯb��{0�P�Q�S�Jx��ƀ����|���4�m�e�V%��ό�j�Geؙ��&��d3�Ful^4�H��V�/n�8�/�r������Y��N�0dB�>���B�Đ�ϓ�kjt(�����|�ְ�o�/��QzDZۍ�s�|�1���ɍ߷��Sm�qkN��^&7`S��hN�p�O,W��S��͵ˎ�
ڪ�D�5���E\�x��,��7�`P��<�"��[5E5�gs��OF]�H��Ԁ�B�Q8c��.v�҂��u/q*,��=W��z�VtѨ�'�L6��n���ٓ�HY^)�}ô��2X�P�y xi6�y\'.���^�� w/0������h�Pm�%Q�c�[Rp���Dz��C3Ιc�v4�с�˜����y��.ŝ��Y c�v9t�)7�-�"��0�ƞ��-ߎ*\�������3��V���J���=	%F��<�Iz5���O@�/ rd������ ��e��RD퇄�m�����I�ԍWid~��"ӋyV�>���mzNs\��"���k�mn�YD�|����<T�����^�Dз�h��	`��o�V��T����DE�C\#;����-��� �Y-e�)W�Ra���q��kD��$���Hc��C�6�Lȶ�&�]�w�gH�7g�`�/����Q��Ɯ
���@qxx�55����v��	��
�1�����hK��f����bvL��X��9�!C���+�����R�Z脹�4Ts�����#��	S�%S<�DQ9�A^��7x5Y<�q	F���O�Nb�ply����,� �7�[K�����M�-%]ƿ3K.X^�c��tq��w��!`�H��]Wj,tTM��9�ߕ��4'��?ז�Lk^�aWW<���x�I�;K#Z���*������w
���n�2��R�B������4۞YHb�sE���/�=�* `�<e���6�9Q4؈�k*�j T;H��ځ=NW���/&.����	c�ۧ>)N�dm�u!�K�=C�wca�|������Z��`*9�F)|[�CC�3�.���ɦ���:Ð��ܴ=W�Zl�
���w�Qk��xvnAA�+�·��6��������Q#m�z~�g����{��bZ�UoS�2A)�
F7}0t$�����:q��>�<k/^��V̲s�a@����e{^x��L<���
,�Uېylz_8����+	q���=C�-��e����A��"�޷��L�d���A��sFa���:�Z��G��X�F����Ȋ�ˍ~���盽.�j��;{��=�}j�%�� ��<��d�6Ez}���؞	��A�>>�� �e���B�o����@zz&h��eCAA;���cf��7�����󏙵f�Pey�9�]�ʍv��@�!��ɉ�t�i��)z�|V(ZJ�G��]ă�I2�[����p�E_��gXG5��k��r
�4;
+��݄t#ָ�@���^��wU�h�9./)�[AB��Nnh����M���>�*���囙���D���E��!�ޔ�ݸ���ΒP�I��Fe�Z�M�SU�Fh���:̕҆F�yԥrL>X�[��x�̲�:����"�������j[c�[o�;ܳ�<B��tR���Ro|�1w�e�+n�]^ 89~ l���Oy��B ���|8]����|h9<��������Rə�/.#��$�R�m�S��*Czs(�]��w��!��&����Tpn�mKA킶�N��
��ѕ��jtZ�g�ؤ�nbr6�k�CxHF���(��bs�q*EhK�(�-yn?P���+��$��ϫ�"���J#���` �AO�/LqB
����d.͆R��$գ}��S���2�H��3�)Q�%ȟ9��_��;�16{����t���i*�W���1�a��$��P�p�B���w�urj�>A~{�dDz<Vu�Gx��_o��-��N[���è|���e��=xN)9i��s�'��?����Z��r(�J*#�6��RW���֨i����-]��g�p�r�{|'%Ta?���3y�~����wUo�?*�$;�c�$`v�%g�y�PoHG4��ϫ��%Jod8�ZS���1��C{�¸l�F�xb�����D�(�u�T˨��X��G�.�����ٍ�bH���l |����Z��꨾��9����޳�oO�凞F��Zx:[vD,!��⺠�Ge�ݶ��s�`v�d��'�h2N���||���YA=�h���P'k��VP�^u��J�+�!��Ln��Q�7�ð�Hͼu�n�Q�����*��jz�SUw���<�T��H'����SD>귍0A�t����Yk2��U�vMK�'���:��NH�j�fY�O�aD��l��Yv���$Ձ>۟P���@1�h}$�`��?��@i��ޝ��#�Q��/+H8�t>�\������~h��=��,��`Ms�<��!�1��8a�|*O�HkTm���Y���	��x� ����A�۟�S��Z���J���M>3�D#�W��9O|	���pe.�������[1ݬ��6�g���^*$3f��݆m��B��ΗA!.�6���<|�`�A�?$�[#��QV��K �g��D�����	ɚ��fX��Ҧ:m(��
�:��`�~�ϱ\+�{�+I~wD݉��xRP�6T
��m���X��\SW]����@�"h��;s�� B������9�Ql���G���!V���a�Q~2S!	����ߌ�]wn�1�}�V�����s�t�����Ԑ%D�c`���ќq�6&znD�386Ն8U���.c��� �MV�Ft��)82#�S�&SK�����{zz��`���^���?VYG��"������e�|�B[���ZG�X��R$ur\`3DYa_��H�'�c����T�����4�ꤌ�����q��f�J��p(�VG����V�a�D�!\�2�����zm�q�=ΰL�p*Ok�վX��h#�;�ET"�/��2F����|n$�z�6����1�X�z{W�n��Z�q)��`�<��&U��*寔	.�_����C�e��RY!�ˏD\B�T��)	�����^uON��pJn}��z�~�k4س��p/�Ꮭ�(��Hħ�B
`�ڣr���%�S�n|+���a�t��.�@Dg�oi���.�S�C�q	"����[�@-�fj�R�XO��iy����-S?5-�6��0�Y{�n�|�9�Z?rv!�J��̢Bƪ6�*�{ϻ���E�`���n�� }�Ճ�J+�w�_�aE�6q0�T҉I��J=�?�03Ƥ�=�#�);8��PE��,�@�2J9e���m��wYqWa|.:�٦�/�ٙϳ�C|����d�S�?:[�C\�������?N�j_��V]s�O���}�q=�i��8Y�j�O�?�%䪊�6��[��l��d��oz��&P��C�A��2ţ�(��Ӊ�sH��!�"�FܢE��W^Xmm4-������4��E�̰�vF�nek�|��voQvЀFE�%��F0�=<��Xe)_I�ݖ�}��W�P�L����X,�"��mC��\�`��#M����>��`1��㒧�k0��P8wj}'P�6(�E: ���@-�� L�����&�8����@լj��dE����XYh�9���j�q"��S��_��4���/�a�v��R�������=�X:�8��s�(��H�>W0��L�R"�^\�ґP
E�D!�?�z?8����@�Y.?��U!���'��"�̛�r�f�<^̋�
���f�7>�̈́�$�-���_��S��BZ$nᎰ<�]P"@2A�	g����&�
��b�E�Z?"���ׅ�_̹�����<ۤ(�>O�Y�`���.c!�Ĉ��q1)��Fd٪w�xk;��*薦��b�Q%�]��dO^:�`&�}��'�HY���#3�u�2ՊcTm�C�,�.���9C�o�W
�����B�Br���h(Ϳ�4M�� bq����s+*���z�e�����g� ��4�-�Qq��;����g�,㞳5/Y�V�oW�S�6�WP*+�/���i�%jP��Ǔ�k�1R�ӳ����7��,n��W�E'���#�ð&s���v�� /��K{.C�>�r&��&HK0��+8��Q	�����8E���x�א��6Q��z7iG������/P���D��>�]��c80�^�W�'#	�F@�3�bnȴ���Z�K��:x>|v��flqd~VF  ��w���-s���{ZqG�kB��<F�_�*"}��0�,����]���������П\ϊ��W<ӡz��L�*�p,)�w���`����,���d���e�*�a?7�B�)�zy�����T��K�ވ΋�!��b��M,�����҉���+?�e0��nYd��Y�`����h*M����2����u�"~�����:㈞��i��̛l�;�E[:-�$�s��}x?��6��)��~ ��\�'Y�U�	? �^�����+�ߍ���5���Ao�Gw���dS*C��$ڙL�����,��8�Q�R�56��)D��]�1���W�b~�����)#t����*�f�y�/����5H�p+DC��9��c���-*��О���{r, �K���g)�RڈUY�洝zU�岊rb�K�����~�������NS��2��p��䓭�kl�|u�
�;�����������Uή��'�(��N��2�H�4�6ԫZ����гY�\3T"_s>K��u�]�y�6����w�C-�mFfU'r5�Bc�j��d��*��p�z�]���m���3���jk�C;\)��	��MC�e)8�oK�0��J��&�p ��p|�tז屇�Mky��� TG��L������;�����Oh���I�'UM��0a�1��� �V�Ef�ڲ9�m�R7��-��n?2ÉNo�U�����T"�y�_����`	=C��a�K���d��sq���|�I�+���?Q}���9���j1#Ƣ�w�0#����AX���6�P
��$QF�����3[�����X3��/9g&d���M<H��TOX��*Tv�a�O�����b��1K҄5, 5m�B�~�Q���TH���h�d�mۂ�Vj;�U��7d��:д[�xR�H�h�&s0����A��ѕ�E�ȱ��(lљF\83���8T���tBk	q��&Z�*�W'd ���*��׸&gM/HWUƐ$�"_ ���� ���<&�E9�����c�J��K�C��e�m�=n	v�Z�\�~�DT.�6'�3|X]=3���ךOj,k�rHa��D���{� )��3�{��%��wm�
��g�>H\�y[�1Tߏ:�Q}�.��
-h���� KV֧�֌�ܵA�qk(�5�`5܈����s�t9�e��dר���洋ݵ�7GOl��g%|���]'�k,��}?��v>����ڬQ=C���(��m� �r���}ܸc=����jj�����m,p͚���V�Є� ^�8v�*�}]:{j��j��/'�V)u1��*��o�H�N��ў9�fP�
�$��hJ����b��7�Lu�x(&Ȱ�)Lf�c?*+@Q�S�Hi�Y1��k5,�CDH�է,�����eOI���h�YBAB8�dfJ�LSL0���O:c����á�O�M�Sgs�l~5�O��%�
(b��V�=}{�3H����8Ψ2���Yl����� �5���>���i��G�)Sk��1�ψ�\wSah���rC�>�y�,����P��+>A��Cq��t�#�9���u/I�E���o=}P�@i�͂��q��#��o7�/�R��ܙ���9rFM3ޚ���ڂ��� I,�qܵV����U���'���l�E`��u���|�N՗o}�q���6��Ktk�`1�>b�Z]�������mj�����'���;DV{�r���ZkӸ�A�?����&�sA���m�,���Nl4��Ĭ�A?��f	=\��$><���>�A�2�� ���j�{�#$"����`364����1q���s=ĕ-0v�
�aհr�>�Z�i9)'=A�y߀ne*!n�dZf�ˋ�0��e���$�nF闙����-V�������%-0b9�|��ؾ���`�h%h%8�j}�Y�a��/Enf�c^����K[����?'�J�%�<�J6����(Nq��Y�ʔ;?��"y`�9��1I�1<��J�C�5�<k�����k��2k.7����ĊH�*�/,�y���?j`�emȕCc�h7S���������L���.��� �xtl�gWQ�!���z�7�����Eb�ƤB��I!]�W~3�^v�h2���pct*���C��&D�DmJ�%+WM��z��z�� w�l��&?�~�p��X�k�`P�4+R���*of��`G_ ��a�c��?�UN� �'��]7{Ǡw�H�&S�pz&(�4-�Z6�/.�~�Ы��-U�f��ķ ��*Qcu;�!�#��\5@��Z@��ۻ[~\���s�l�/!&���Fd��)���na/�V[��njr���TQg�N}3���Jn��5����#On---p>�Taw�xI���u�⤐�g�T
���@z��4���Dc����t��b���61K�0�j�}-^�Р�ѥ�g��,�V;�bb��f�����[����\(L��V��� ��F�AѼ�.���v��q��g�DzP3%�����'���������nkL������&���Wz�Y)�w6Fr�l\��g����1�tO[~���س���o=�h��͖Lȣ
�c���۰	�H�gY�Sl�/<'��.��:��3����{��A�Ʉ^�"Nq]ERF�#z�T���R�b��ݴ[�d�|�L���ݐ��_҈�HW������ޠ�/��[��Ҩ�}���Yb�~m��#q�ݤ��dA�����A��ʧ�ֈ�?�j�h�t8���ۄVm��zΧ*gぼ>��³�r��SQ<I٤M<K�d�V4��R$�������A+�����f�by�b0�57�=��
����űQ4�^�����J�$T��X� �s����m�'�Z�i�2h��b2:ν���;`{���X�P��7�qZ������vu�h���lMQ��g�}��W����k�K���L��B���d�	U�!a�	@1�,e��D��t�/���^�+d�ٖ(8}`����e�v���pe�1�����p��]������a������`�9ǉ�����(oq�ܞM���I�b"+��mG0�U(�jD�m(�w�-�U/��#�W�/RU^�ա�	Dv����3��&�y�s�}�o*�O�f��N5�^�s��9]���w�!�v5���T�Z7�:ʓXW�i�,�o�t6��SzN��gmQJ�a^/�Z�KD�BB�X1J��~�
*���p���Bѧ23��3����2�L6&$j�\(���}ֈI�f��{8��������: t���Å�ܨ�M��.�jc�`B�h�>Dg%��	cW�}ii���9���L�U�m�
G��v��O�Sظ$ZNA0'�]RXH���?F��f*	���򆱎�����b�.=��YeĻ�
��Z����ݝ�qy ��`��\�9`z|��b�;��:@����r����,J.�m ��:A�0����XH������
so� �W�`�A\��YG\����s�U9�p�)��g�����0X6�S2oQ�#�����G�-�Y/�"������_5��9J+xs�>�1��)��?H�:t9�Ǡ�1:�$�(7�Y�dK����Ҥ,B���+U�9�r��� j��W�l�uu9'rx����j��� �?9�E������s�ќZZA�z��-�_��Q+�|��,'��%}!���h襎��@�=� ��U��e�e����\��q�Η��S(Ҡ�u�����v�m����*N.��0�2� ��T
�T����� OyV3�s��v�spF�@�g�MV-'�2�iU���QQ��˰�3�
�T�����δs�3�\��[-��Js:zZ6���ϔ�~�z�6�n���SowɄ�lYR�lG��CwW�6�i�vVI$�1T���3-z�7"u�t4q��(�=���%�xU�}����G�՞T�:8��Q4
V�?<��^�l���ֽӀ󉆱>�BKg,? ���ν�N�d�̒�&6�aY�n��"���%��@�����#�����˨��9���*B|(�]�U^��� ��V���e��oZ!=gj/�v4�T����JGp<"L�yb5(w�ME�6���I@L>&nK��˲�\6�/���u>���,�\�9K�����2Z#Dl/���Z��QfHx���J�ث�J�IsJ�4h�I�0|4�5�v+X[�S�.�v�i��	['���lsuK�����>�K�M`/�}�l�믛��ͩXB�,;��=ڊ���^t���( ���`�2B�aFS���<<���V矮>戞�&��ڧGg�{�
ƂZ.�����b�����2��s��I�q�����)w8����7+�\WX�������^1���!��0��\Nd��a;t]7�V4�(�*�N��m�9�FJu�Я�K�#f������<#�u�$7`�U�����$���}%�W��C����n��L5B&xV�s|q�;Gy���6�ǲ��k+е����C����ͦ�I7Ѡ�CxQ(�e!n�nDNkqX��`ryC'2;t��T;3U1zE���L����Ԩ��ԥ��wy)�C����]T�	v�S�U{�6X�s��5�a��v݋������]��-�α�$��!��t���̝E+:,d�=y\�m4��X�eX�1K����B鈈qk'-�9��/���E��.V!!�&	��S�V^��[$G�@TÊ�d���j�wH�Y��D��ɗ������ԞW�^BdUg���ʰ�g1�˼���`?1���������X��G�2R�-���1#���\�*�eXHښ��">H�BX~LaM��`f.��j����)��:�Y��|���+��ٟAR�c�k8���\<N
%r��i��rƻ� ��Ǣp\�
�{ƺ�}���1�o�rz���om�B��P��
n���7�&���q_b\���2'w��Xx��ux�hT3
�F�]tX�yUceY	I�Қ1 ����~� A�����<�H]~��o/=�?�I��Gu��:�V��>�Re���mr��pKs��I!DR(<#~�R�=���_�"���z8��D�3�˓^�k)¾�n���nPW,l�TY̖(g�g��)�8/�I��Zs��i��s/���uq�T%��cN�����hk^����b�wM�H
tB��q.���G�30lzg�b�K�*��J�3^&"d)д@|nX?]���e2����Ī5̹D��5YH����@T�5���ɸ��v�mWl���ψ��8�^N�Z�
��{O���uȿ���ȝ���c��a���zS��64y�i���R�Ά��T��(B�C/�t�(8U-u�c[	E�c�Q7�|yĲ��[����ʫ�:@��:ۏ[h��K�����l��+c����@�K(uz�������?����i.� ����1�.R�(S-p�{�L�L9��WwO%��7,����>a]D��{{�Ў\�2���&���'�N-����� 4�n�-���z��nv|�t��.�&ٱ0ٽB���2�0��{�d(���UY.я�;�j[���G`=ljA�Ri�X����ƀ��w��N�{���y�Sj��jM�h�zi�_�6.κ��p.�f�ɨ���>+�p�c0-8���h�������^ܶ�j'�7X�:F����(�/K콠VN�s�A��
�]�ݼ�T�D�`��B�qLnP��&
uꦙ�����a�y�h.��ko�g�e|v}��Ϟ8x��@�q7 Os0�^i�z/0fе� �͛��%B�FΩ��ˤ�	��������[U��v��ɷ+g�;�&[���Q�[�ׅƉ���ɎE��*��7" ^���VP���C��?󭱻�#90����N����z�����S���m�,��+4]�sP���.�V�Ħ:��G�7�~�:�=�0u�Q����U{+%n��F:��k �A�۔�ѵ���@)cv6;�f��D�~����RȲ]2������_J.�~����]&��;H:�5�����T���9l7������Ej���#��  KL�:�r0�i��`�ep�J'�r�������rkˡ���$���G�N� �rI�Op�Vn���� ��� �zЯ!�9C���Q��#w�q؋@UOt�s��X ����Ϛ_��b�U2_PT�8%����]��@���E�r0�������CPoy$�e���¬5�5��[�R�׈f�B�1�,=�c��?��YK��緈ԍ��^C�n�rU4�IE����P=&���l�Ǎ��J�W�x�W�»���=��Ղ���Ư:�ݘ��ܝ*K���\�R��[i��Rzf��=��c;���,<ʀ�9	�8�0��Nt�:�a�����;����\?�ŀ�WҌ�`���?6���h��S��c�'zsި��XJ��us���u����EJk*[ ����v�z��T0��/נ��G��#l����]�N�����~_�!h�j�(F��!c0E7��$�wy���(�W��%�"�ň��4`7����͙F�a	n2�O�B������C|6�y������*���>Tb�;��e���O�	�P�O��3>�؅a�0�GG�rI��͇U��&�u~��S�7�J]b �&8<�|���tfy�_�v�M"�j�?����N��B�=�g q�hX�8���ݺsܴ탸a�+�mE�*¨-s�"��4�u���8�匃�}0��|I���`%,ƹ]��n\��/���C�YŦ����\�
Kt�z�,$�����vr
�[JP��|�="� E��a���J�&9�d#9 ���P�%3��6���\���(4��;j�;�K[ :)Ua�l0��FRٖ�ݹ�zY_�.��+cf�Wx�����_�\�{����Ĉq��g����C%����@�v�Uh�0Si����^�ԶʂvpC�d��%��t��[xH�p4�A���GO˄N5F'/��fC �2x�rVrʄ����1K����z-ŕ	j�&��*BP�S�i;�g3j�F����(�J����>�9��<]$�U�֔�)W`��T��Y&T]����A��1^�P�ϩ),��L6E>C;�ο� V��4�
���RΫS�<G~��	eJN��r����u�e�-�ȱ����HtШ�n�ν�_��$���<�U�#O��V����Cј��X�s�K�|�B�/�A���d���A����Iv�*t����x��/fǈ���V7}<��L���f��ѡ��R�	��b?-�C%.@�[�;�ݤ�6��o����H�ֿ[�7W���@ρ'."]ME���g��;��E�W'4�4�.���S٫�TQ˷����;��X���`2��&Ŷ$��z�ûg��[g�!4; U+ֻ�`��g���&�-?�tJӊ\�m r��r�1"y+��n��ɣ��+<���G�.Q�f�$�d���Y�JM��M���GlRo����7/�B_� I|v9�Ha�6J�(���<��7v�ak����H5L�DĲ^�~��޷�6V���}z��?�X��3�����&���ɰk��{3B
�kZ���*�<�}���K(���P=f����[�sV�� �U�ӂG��7|=ub8y�M+Ϭ����^�:/�����y�A��V�re10�ɴ3�P3%�L����e���m��Ծ���ϻ�-�WOC�E�©.S�i*�f��fgJ����ĺ���)
VH
$���r[�]6�.��*��X�m��A��������޻���k�@�ϯ:ΑlՇ�a�?�V���M}/e2����(��w;1�b�v~ζ���)�g�_v�4�h�+b?Sv�!���M�p������h�[U�,�}�$�\�� V��-�[�ǰ{�̛�Ygv�O}��Ը@��c��(�%��oBS�騚�`�pM)g���9pr��Z`T�5�tp@ֺ�v�alz��g��U�����m�|�	+�,'����ha�[fc7N�+��-�n"�*),"���	��	w��_���}T�N���[���oyM�9�žG:�c�F�MS����=���
j`��`ߜ;w��<0r�>��!f|V������=:r���:Hfd�� �b��m�!���B�`�'4�>���V��	y����<�W�ר4���Z F��L;o���F���:���a��˼�r�'/$�����9;�	ʸ�'�L�} ��yxWd.����!v��1���U���� �:L^�s4���~^$�H� BN��hWy41�ꏩB�Az�ߕ���Ү�uJ�ySd���6�o̴R�ɀ[���Y�o��^����j��.����;�70_ލ@���S��v}��B+��j�M�z�Õ��Y��4� t�1�_���3<��}7��NhKo�^��lasf�s������:+�\��`	ZУ�g�a:����	�z��>I/H���4R_|KN��7�����h��R&\Ƌ݁��BW��p4�K��n�a�|l{�CS��d��uY�1�"��\�Wu�
W��Ry}��	����J#w�=F��I��M���t`��D��C����8��A�n~�?V�p2��C���f5����X�����3�@ŉ�W���J�o�cd蕻VW�2��K�XG�̟+�k���޶��Wv_�v�y��|����b�OT����2�d�q q���*���Oj������'��槮MJ*�hB�#m��� ��������y�����V��2�?X���=V
isb[<�6�|���T51a��D�Y����Q��Ok4���r�e��IƂY�H�99Ѫ�Ov�p�M0[ ~�T��u�m^�ǃt�toj�-�`�n?8|�dE0��kiWBz(���R��]���!m^U���P�1)��Shy��2�%��fty���9�i�?�k��ֈ~6�n��CN*��Y3�h�5���'���_�dС�:���v/⪸*�2����;�F��R�%�;���r[�6@�^GS���$�8�3���B��G+�P3��劼�r�'ps��I�~��)) ��d�������0�D�N�LC�8��Vu7l��` �m���ܡؑ#ۀ�y��d�`�Ɓn�n��`t�O᐀��'��%�Xg�t��\����P*����:xĆ-d�\�Ah@�P۾���\x�t!�[K���-j���hlV��H��q^�����,Eo��vs��w�.��Cﮓ���ɹ���9#�����Q?�}���Z7��J���\���+݈�zE(�+��~���r�9�m�AmVU,���i�&Yr8΃6��-��C.<��Ӱ�����S������ �6�[�MeG�;i4� / .%��yKbk6}���������y'zIB��<�x����~$��i�)Y���Sa"F��l�:A̼�I����<���̙�dH׵�Lm˜�=�g���.���ss�gT�* 7�KM&�=0���;�%0U_ yy�AT�tQ�ڻ�%���
�6��OAV}A�@��Xz�ʂ��0�n�6����`�׆�D��j�=�����=B�&��݊n����&;�?���&�MN�	�O	,~�
���d�R�{���`��J����1w0��?,���?��`S�H�/�d��{�i�A�=����%���t[-g]�+��O9�\�oA�0�&7���%�Sa��wք��GH :�^VȄ��.4��ޅ/��T%s�;�,�S�e�(ۗ����.Z����M�!e�p�9r���&s�x}�#aP~�'1�C(G���_��t1��W�����8��9�N�o�K��A=�Fצք�]��cH3�c���G�Ƹ�\�쭃�p������s���Τ���r0T�i��!1.���ho���'M>��w���z��4w���0��n��6��eK�rr�ӚGa�p�@�����O�8ѳ�;����,�z�H��>>�)�W�Lw����v��hU�p!�U"���^
���z��aw܆�wf)�C�H{#�b��	A�"^_j6�Y#�K�2����qӧ �<_BR6¼��<y����tj��xƗc�>��{�*���!x��g��������?����sRw�b�r��$v#�\�-:���P����y�a�*�G3G��jm�M�:p?��F�,�b�5~�Q�?������N��_������7w��^���-�ǚ��c��Q��"�b�*^Fw�9}m��,3�a��Ӷډ�cP�y}Px��r\ �)�9t�o�Ā2S�\�)��<���T
E��{. ����>�����i��,�kX&�)�h����M�SjXL��[���@=V�O�}�m���T�����_h��VT4�j��ދ\cw�<�G�>	��ǯ ��Ɔ 7y�8ZӴ�i�>�CF�'�'�M�%�/�� ��I%�+oU�0� ��}��HF�-px&q�"M���Z2�rk�O0z����_e�ki�屮@ $mk�$��S�YkBq�$�x�l�CF��cN�����U"h�$�Ւ����ix��=���o`-�6}2�>�K��Gy�tīþnߒ�G';�;0e��E�Kh�}�/w}��W�f˂���k��	�YI/����w�9�ƪ`��4�Z�/cXǭ[�iN*�*����s�1XBL��^C ����%-J�D�6d����Ex�^�w�k�	H����%�)ۢ�a�r��G�D b.�����q���������8y��q>�̂��z�
v��X�k��t�v�%��?:�Ml������ߋ,�=�S��#���(1(�ϔ��C�M�%��6��\���'��S����0��J��4W�"�)H�i��)s� W�
JU��ە`�4���D�1W��Y�VW��z5�^��o��O�X~�>�g���<>l�^L������H�P�z��H����B�s��p{�b�Q��{�o���!�:!����SvQ�	�;㊞�E�b=>��wq��l���p���y��/߿�=L:x�:�zr����E��s�Kv8�gӃ���sE�@��z�[�c W�au�W��i��h��9$�̊b��E��l�|�D�M�9��*o�&��_$;��{~g`pΐ�@�־L�T��cIr0hJc����nGL������]`7?���{br�ڱ��v���7��s��w����/h�`�wzw)����W��?~�G;����;IKl�C�n~v�r���*�M� is׍»ට;^ E�1�o!�򓑭���SWJf1�cbR�d��;���V��|��H1�:¢�G.u��l�w�RC�S��pn�q\��;Y�R�p�
�\_��VzH��s����kT�a�xq.q�,��f�[1gXy@L�"���R�Q(q�-�t�u3k �\S��$�:��g�fZ������wb��[�`�����-�5M b��՜�u{.&S��_�F������oD��S�)�]ׂ����}�}<�P���IN�b}=�ɤa�dL�O�_�V��(�I�Fq��S��h��ZA�+ei��;���g�{4�QQB'Y��,�Z۬�=�<���;��-�oh�r4�"䓺v2�T���l�2�L����b޸F/t�e��F	���m���yhi�Ì��L�>�1�8|Ʀ�^���Ȝ����Vk�+��-J�r�Q����$"�0=��T���ǚ:���F�������TT��h�S��7'�:]^��op�)Yywvq�zv������^j(�_`�A8��(�8=�61q�{a���76�И(�*�C0%�.���x�}�J�M]X�{z?s3��!��6�x�٩��;Ì�����i; A�R�ܽ���Y\Q��1j��D�/�5@Xb���^�$%����ۃ��	%;���ެ�}l:����aƳy��ٹӕ�ɧ�+ȺB�f��M$�U�|�}g�Կ@��/��9	�v���S��@-/�����NC>We�)�q.Q�5��qs�^��н�s��k5$��[,PԹ�kq�І<R;�Ω$="
u���T���Fk�j�Ek~D�I�_v�L�}��9Xdu�������A����`�eH���޵g��23>8J�����y����q�QQMVn��(S�͂��.�����-ѫ�b��x� �mß\]�n|[1�D2<�6
�p���'�ǕT�S�m�#
��A��Q �` �9�<&��
�n)d-�|
�o�i{E����!���|��Bgiy����(� k}8�	���V��M����Mp'@���љ�&(|/r��O������S$���x��;����=����R����'(Co�BcA݊����F�5����)PK?b���
`���_#�D�J<�ç����H���#�" �☲~��O$��?��9A�2Z�>���+*�6����%������f���� �=� ��1�>"�f d �O�f�z@�bC��!�������Av[�"p�H�\�Aq�� 4��"�67A�Ð�	.�üF�ŇSS�����<Έ(Ւ̐m'~���0%"ՃegU��)���_&T����&J��?��+ը���+9���.��K@�9�ǔI�D�E�5�k��5j\�w���v�i�k�㰏0�a�m�9�P��d�����C�T,~���E?1����4M���mS�x2��C�)g��gd�,�\�w�b�̴��k@��w�����k���BfBw5{r(lKcD1�0�,�U�x�vR�:	�/��`Ks_�>>Kz���� �iU}�m�^�[K2�3hԐ��Q��.7�!��{�œ.{���\P,���T�S9
4��P�غY�~ �eC�K7A${	;.AZy�t3�����xvF�qU� j�h�'`�ym]��Gb�.�K�>XP8��%��
�k2G��S�:���J���s�!ZH�U��`l
Ǡ�y��iuI���6f&�Da����gj�����S ��ŵ�/<^���NvJ���i�#��5?Kg��X���e�ɱ��/aj�/�yB�1�z����)�q�EÛ9���zV��3������&-u\�h�9c;�go���%cVr���E�u֩C�&Ů_܀�D`l�Wi75C�����%=�_>1!;+�qzI<�j�;$uA�����O	����F��@-�S�3Z70oV�!�y"N�Hj�y@`؊��3��HN��=��!P��.I>��՛!�]@B`�8�Є�ӏ�R:y���7mf)*/I�����uw43���r�}��@Y���*�&��rq6��>��5�wvZҒ�x�n�>޳[�JR
	B��Q'��:jU��#a��d����Z6~b�.��C*� �)��Rယ��:U	p�~��$ݸ�}����ڼ�#�ZĆ��m��RГG�eZ�??n�>���O�����վ/6����&��懞r�!���d0ʼY�/t�:XǤ�v�u7����>EUľ>\|��� �3�K)����Z���4��'d�T�F̮]-�ϩ��3�%��ImJyz���Q��Lͣ��<�^A�C܇	ԅ,GJʤ�ǥg����ۊ��5�͉,�Xhv����nT����	s���N�u7�����A~���#^`�%:*��k�ڊk���{�8�Ya*����O�l�m4��QhR�mf�׿4X��`���,.��y� 1�R�@U2|��i̋���(�@7MC7�?j��$�zS���8އyHfh�.�NK�cƠ`�2Ԓn}��~oO�W锉�Y@�!��6S�K�9v��t�
��B)�y����aA���p�&N)�8#G�0b��C��̩y9�:���mw~��./�4.J��I�}f�=X�#��O�C���Y�ss�V���"�T��ʲ�w�k蜌��M'�.�/b�p­�%j4�6K�� �P��G�苐OkfI�6d?Z�*�y+j�"Mh��UC�%���Y���ܢ<��e)wYkg��͌yaZ y���tb9ɒ�#<ڃ���Pǃ$�K�b�2t�}��ü��|��*>4iKi���ڛ�s�tÁMk��C���'�*�	�����?s�z��wnv|=��5����c�Pfug��;f���x�<����!Д��䚬�K��R'�H3W���&p%�C�noe���%5V�y�@)X����>l̔����-ϨM����R��%m뫿ů��W��I�//�I.^�>��Pn<��[*�V�s]��5�k&����lR��	�%SȺ�ZGI�TZfx�M������~m�x��r�Q��+P��Kgy��9���4V-72�-�i*���L+BIU���[��N�����p���@�Z	�a�G[�Z,YP�ee����Ģ��4<������&.�U��+c�ȕN�&���@u;f��Qe�ѱ�o��BK��-�CIҍG|�J�WK�X'p��s�k��SUy�sy#�v���K����]�����՜�W��w�y&x��y +q�.���yh}��[s�{��c1tlmS9�[��g��絨V�"n����U�`��������w8ż���<Q3a��X6�MZl�MsJ�*T-2�,�n�z��E�8���G��UHX1Q���u�`�~ޛ()G�#�b؍f��0���_�)�41nVжԊ��f���F�H�k���> ��KVL��V�z�+���#D�m}t"| �f73U2%��P`~|��mf�J�IA�FF��ɽ�[��#���Y���l�d���	�P��} ^컣n���+�kލ��������G��K��Ԕ �Z��UA�3��d���]+`��e����߼�p#��,��_�X�7Ep ���/��K�DX��2�%
�2���%!%��|m�O
��i^�Z4�D4�~��g�MǇ5�U�F}��7)~wb�<�~ac= ��[���4i�d�C�� ���g�,4ʽl�\�4�H�!~Z���2�|��Df�3��g�y��羚ZS:27����W����jg?��4<ԩt�Ӎ���6��O�������x�3tT���H+Ƞ
�hTdx���~�o�3K�9��C��R����0�]	�&��Fzǻ����7��\u�k p���PT�����3��|�têZ�w�3��V�\8�y���
���P.�b�e7�`Z�v��υk,h&�QQ7���!+�|#Β��ј
�e#���_;ن�J�d�y����p?*���F��Ȱ��|�jmueS1M���=����/��oC������,�����o���5��-����?���8l`�+Ӗ���C�l+�k��2eG� ;���T��bFG��`���R	�bEͩ�l��_+'=QL�����J�| ���1�+Yǆ�gh��Z�~Yc@g��OU;�t�ҋ5����*�?�t'5V��N�V�������U�|<wʆrxK�O�Iꞵ36��� ��p'u�8ƶb�͞)D���W�q?V,�$�!:Ϊ�)��zxH���z����W��M> ]��@.}�߶w�aP)r'���Ue���4E��?@9��\��(��9�9qN5�����H+��O����S��5?�E�"m�FE�6�I�S�Vh�}��_�# �s����"v��:�V{H���Z��irAowٜ��H8ޝR3�/����%��f#njy�
E��D���Z8�����!M/��r�wʿ��]�E���6��35/d�:/�@���ђ�C	�F�TR2'���lw `��'V �"w��Y#~�x�ͫeoeމ��b�H���6����S+SE�&O�xON`4��5 �x1Lo���i�á��u2)����fO�I��ד�����q�Ta Ӥ�i���^8��L�2�������
���S�t�zrGX�y$6a���O����A�|���91/eM[�����t��x ��) �)G�~�/<μ�M�\춑��'�L�q>a�.�M$���S"B��Mx �N�%;AcF�n�=�f�rsǭ�n/j�a��6x7���()R"I��a�>�f��X�5������Z��S�P*���;��5C��$������d�*~�N5g��(f��&��%����9ڗ�M�"�y�(sv�H�l��Orn-�F�f�bun޵!@\H�� p�8#ɕJF~9n�����ݏ*�Vx)-��-%�~4]��#}���ϳVY��H����������kNj0�˻ʘ!�;�=�h�����q�"4�y��qM[a?�%f�eJ'�5¿A�ܤ����~���9���ĝ�\�=F�
K��	��#'�^��(�d��]/K+
8��I�Į6#��O��~��l%0T��§Uꌶpb�a�|����J�mK$�^-��V�J����2ԕ/�`wϿq���e�x:a�<�6*�N�k���>oGŖnK4-rd��qfd��� L�ne�u��2>�Kh�,�Q,�]Vl���c����S)@���^4�2 ��< v�Z�r���N�N��X1��A����r�w�ΰ8�	"p�~8�Z+����1ǋ�5��u�痑𵞒/�V*�އ�޾clʊС|��VJ8�ylL�[�i������"',h{�aʶ�Y >:���:�la�C{�5WAws�֔���sF��m~�e5�A҈ܟ�耙��`^?�R�	�K����#Z='m��˚^?��:w�O,��kҒrVYy���ؽ�;D��َ�p@�{�/�P�#����R-q��ѪS��*>��W�,#��5 �|�s�ֿ�`���L�Ag����x�jz9�kh�
Ӳ
F�*��l:��!�u��N�+a7�[�b����7� vhd3H]L?>vu��6��V�ʾD�J`��]������<ݚO�{�����`���ZC�[�Ӛ�үo�˷�^��u��]�&Bv��!l�w�,���C)�GH�Oq����u^L�p�q�.�c��%�)p&�y�(�#�.�md�Q����GQ@��N������b��v�)�Mv�����h��
���������s"a����ޭ}�b�U��bɍ��>�!�k����L��~j*��:�6ú��d�j�_N+�ȜsU�@�D��nb��@���A#I�}x�5E�$\�@��EQ�2���_l��驤���ݱS���O�&�L-����˛����U�:��d�
����W|�ߟ�El��=״L��0g��ꋓƢ�"�
+�e�ͬ�Љlc3�8+$��Y�� j�߇0jF���j]���{��J���W��:�6�_�ǃO��j���궹Y}UШj�WK�Xn�_�^�QI|�J%wU�U#�a�dF���!(�սP ec�"��r��<�0��.��](t��/�6���1zǠ��4c��4�D�}\�6\���M�3���g���ϕ�-�J�jYJS�Q�{���a�9�J�x��q^:{p���F.�`�4dƛC�T�^B�P8]H�o�&��[��!h忲O�v����d��%�|t�]w���>���!�r_�#'�b�]tܡk-7	�Cvp7,f��^Fi۽Ⱦ�]�6o/�
S��L7�E��e�Wv���l����̉߅��<JP���&�	��Zj�X��a�>��ůY��)���2�5ֺ'��WX1����1}��6���1pr^u��>0�GX{���L��-�wK��2.L^�w��3������(C?5��1�@g����QYG>=�<H����N{�1D�������y�_־�7�]�JrC�(��;>`f�l��j��
Nj6�NBEX�;}b��P�<��_�RPGL��� �ۛ��󧽕c)�:Nv8��N���d�G1,fn�m�)�5n�$b?�����U=�z��Z�C����d��i�'B��WT����#k>�kt�F9NHg:������кI�6���C��,Z'��>tu�fs�׻�RhOn��ݬT��Rw$e�Y~�E�^����n~n_B��!������I�z�\h8m���N�m���K?�SG{�~�����nY0��fL%"<�\3K?\y�/�LҒ77�mvHN'��E@
�}mu�4o�M��ӏi>��k�W���Jc�m+Mz��s�;O�K�����39�կqvIA�r>�p&�q�H���8e��}"`�U� �m@r�	B��Θ4Ȓ������z������"������k.��s{�v����M�#p�"��w����`����݈\t��*�\IOV��Bj~Y�PK�U��%^qڢaE�� ?��D�-�5��_�d|���9�:��(������;�x���Zzt�f|?%�|������Cpf�F�@����r!^C�G��N��h�\5.	��(�~��,c�}GV�����_I;����1F,G+��?�m�ܐ�ݿ�������-n�-�q�i������>\��F5�
$/��t��-OڌYS�B:c��K�']�G�Ӕ .k�&/��]SR�ρ_��m��j1�F+�؛-w��<�r������(� *d�U���L̩aϑ�J�̐c�1Z^��By��V� T��=�8.Q��mˇܮ���Y�
��v<#��^�~ �����;f�K.= ��}��m�����Ϯ�vE��(7
�$,�둏�@�\5����*��#	�u��
/�!��(��u	���@�Υ���N�#�=�_F��wuU��8u[.�,�A����2���O�!��#@�a��a�Hn�{�ܪں�O��?�LǸ�$_ x߮�v)Z�0͗�"�&�yN�P��3p#*q�W��#�)�f����<)+BB�����ƍ�Gً��z���Dm�vHD��֝��p�[2�EB)z�O:eX���	�pؕChg/g�����$∓o�VN���[�e���2d,���	-��Y�ՇխM#�۫�k�:�K!�U��˿�-�a	w�t'���N��}܈Pag��MVoI_��y�3ςi[5�"����,N�s����.�Ī�b�dnN��=���v��)��I��xK���.jc���4i*wM�����z�!��:62�&B�ҋ&�7'H<g�)�K�Β۾v;)_��jR���܌��q��u�P�qe-����W�Xn�l~��@���8��d"���*%�nO�7)B���LB��i���A�FỒ2:TXpW1����m�ݯ�����]��z�f�krM�g�b�4�@I�O����S��?�Ǚ��#V{L҆�{���\� ������g&H�n*Ǹ����*w�eD�����~+@�r�	|v���^�ď�E7���C� ���^ê�)�9J��!D�n~��q,jf<�h�g�ҹw|�\w��V�,��g����ӻ�Pn��(<0�(�/@�����EQ�y�hƀ�. 3c�m���^k@���XY��)P�� ��iT۱�e!��*�q����o��)-�٧Ǯy2k&L�V�O(*[����bS�*�|��o�\�%$�<{��"�-G�r�#��E��ې���^��㑣|il�������cr�U�ۃ��K�H��3�2W+޵gv��j�0J�G�z��yvW��d;Ա�3�J����=Z?F�B��Wjd��p��! �>�U�<�Ԋ�B��v����A��+ݓ�q��TDuE���j'bq�{����+����>-�Y�Ms�c#NQJM��N����J�UY"��f����j ��!�5N#��~�D�=Ƣ5�� w:��IL��E#K3�k�G�+h����w
�c�`�F�"�`Ȩ=e�~�wp0`�{o�.�NP��t9	���.��!)�2���}OǞ���&���5�� /1`�T*Ŀ��?9�U�#��-��Zk�A߻���Y.����1��e,��2��M��P#Ͳ���3�n�>��џ��\�g�["�yo���Vn�$Y�)���5�r���%?:7��Ia����[Qj�L��&GN���C���/��k�±!hxn�϶Їx�3 ���B�ւᕮ4��Q�f�9z�zq���^��%x��6�� v���w�^�g�m@�ٞ�c��� ?��a�T����jk|[�r�rݙ�/�Ul/K��D�a9���l?�N:#:�4M��3�wj�8�}��=��+!<���~�Lx�����R7HsC5K_hJrd�u!MyW�x�!�����a�.�T[sۨx����j-*��D+FS��]�%y��A�Fk��<���RtwF�o���kk��7����V�k���$�,�8c��G��W�L���K�.U��A^S�ˇ,Lq�:L^S�Z�ķ�
�$m)��h"�����5��3��So��I���m��%��.�V3c�����[� {�=eE#Z�" z�eO��Ǐ[<`�IΕ(hb/u��_}��F1�J��)d�g�N�B���	P,ӆƬ��(-��qE/�F��a�d�I3�U_Y�h����E���+����
r^�K���Vw�\v�x�r��zs �+~�y��w�y��΁����6��Ky[ń�������?�Hq�e97�T��7�����J�����BR�ߘ��Z���Z�`D�;RRZn+M��ҹ����kԺ������ �=�I�:��C�np%--��M�ՃxǓ����L��p�(�T�MY�E�=��	�&&��� ,$��.��1��>�K Jy���o\;�k��m���!��phU��4#a]'ȀvG�/����v�p�:K檰}&�6t�2Uh�V},l��ɸ�Y刹^J� jC:�:TQ���W����!b�����r����'�ϵ�ۺ�]lg�9jg8~>8��n{n����v���)�tu��珃�w�����啉M��1d�a��hM��F�^M�tv�oH�R6a]�L�iڥm=�f�@��ń�5�AxR��D&TA�pnmp;�9�q#���麶c�s�#z��(�K,f��c�ą�{�呪�u,	�����Q��xm�K?Ї�h���]J�~�dQ��b��l��=7�s�Ʒ��s�����!�T�,���	�A��f��1U�Rf�e$�3����>rrvl���B#�l��#o{f�EN|C�OQ�x�;�ku|���u `�U�위�%�R/Git�f녲���@�4��Ll��]��&�wQ.�ZF�F�L���hL��t�TF�&hp��T°�>t�����E{�]�����`�K�U�v'}�"�,6��}�5?�vܛ�gE۝�����[�Y��~�B�+�)X��X��]	��Lh��-:�8( r��M[W>��0�ʥ�cN*�魥�ǟ3@U�\b��)��)&l�lf\=Zo��ڇc����I:�N���T�������P����t�� �5J�?֌rk��Jg����u{s5��I��{bD)�U��C��O��Ͱ���à��>(K[3�C6�CE,�~,��`�po�891��BpMǣ�su�*�/�PG�N$R����$Ց:¾��'w!)]��F� G�l�[N�iM=�. @��/2/�O$�S�o�ɽ�=�O-��m��o��Ӆ;��G
���9��#0d͛a�����B��*�����F���3��>��!��0�W��:Tb���T��Ųz.��!AlԿkK�(
n���d���8qWʹ3��j����77&�X�f���I�`�$�f
>�[��M3�i/��a>/���K�O竪ez3��.P��V'��}1={�\5��j�t�K�
�����W����	�\Ch�bK�K���W��W�D mR��!��
�����~� @[�p�=�oܽtn��'3I:g��쏝_��(�4 =J[�P���E��WK�>�nc*�]j�'�W�S��*��H�@&����-�K��E؍�vV�����Q!�!;��+a������2���|��.���E��I�]
�b�E��0��hi+̖T��?�y(����f|� �AEdqu���}I�=I8|����]�����K��$��	4'�-/[�57�U�NY�l,*��[���R湃(y���s�;�W��r�Ԁ×�����AS��kxvp�<��F�����}M~o��.!5^�Ńa������O)
�%F����`�к��Li2N�/8M���EP�h<�_���J�K�����\��� �����!�XsXo���n2-�3����a�aҹ����4H�%��1��g�4�\J�oF�q2}�����qH�_�]�~:	p+&^0;OJn���r�6���  �d��n�E���F���v(k��t�(תu㦺�L zrJ�=��Ô���շ�=Ur���F/6c�Ρ���F|�Q���n�4&�=�����/�?��j�>n�z��Mm�Z�t�[	F��*6���#)~'��ᾫ!�K����%�����1q[�լ�r#�
�O�{P�P0�0���r�A�B��Ot� uU)�)�8�LR�wG(�����9cH���FJNY�4�Z_`�s�u ��ol}mL
US�na	l��Q�ޱ.�oB��t�Y���'1>�9,&K�&��/k���6|+�AQUZ�����o�hWM+{Hu��Q��?9�9�3�NO{��T�7�$,G
A//M٫C�7��;-���\�S��: L��͔�D �$c�㊘�U'ah5�� �h��,�O��"�����f� ��x�ګz|���$�����Y�g��r�3P6�� �Ҹ�r���B���>��ݬU&`en�@�ܽ[ȓ��xS|
x�4�xy�9�p S�Y]S�����ɖ�[2����l�A�[経�Hd�'��MIk��b��h߶e����9��#|[����܅-Th��W|)����PmP�fފ+�%��E��r�E���A��2C%3��%��y�e���T���.mߚC��Z+JP��,�n3�0�"�����r&�/O�-�_��+�0���|�����ae<��O*�6a���I�dD��j7��s �4�h��j���w�E� ��TɡG:�������\�F�s�,��(�
�/�#�����v�y�#�'�G9)����m��^�%�8���"��j�
�-�iH�J��;I�x�'��)�%4��+���d~��6�{�J`�~�����wT�?^��1D�5}O*�A�rL�{o.��5�R��FL��8�����y��`�q ̤����DŹ��y���nږ�������\�L�Y]Sj�.��ƨ/�g�)"I@4�n߯J��pPY�)a$��;'IyLك_�9b,��8*�=o�n�h]_�ۜ�����.AɆm��tE^��R�����	3�^B�c�S�Avݘ��_�@ܸ3���8[.���e`6%��㵬Wz�X���&��(�A�ڨ�&���[���@a�,X�_h`��p<d�9b�Ʀ�?t,4�Կa�#K��:�U0.�Q\.�77��o��ܭ��GΠӬ`Iȍ��=�\��ݍ���z��|y��O.��\�c��鮫�Cӑ���2�HAr��FqUW���(1�l,��gqS,ٞ0π�A��͋;Y
I���F�U}����_P��98�g�r},�}]c��06��N_��m���WӘmd����x��A����w���:k��3�}��(��^��U�F?_H�
���k�کW5﨓 ��2��@��l�@��o�ɠ���?P�4 ����foKq�fM�.)�4Q}�n�D�J�.vj]	���O0קh�k�Q��w��?8h���5ٹd/>-���0�NQ��!0Ɇ� Ӝy��d�X��ʦ��5�[?�����%�@[C2��J�4^�>`�Z�;k� <����@��ޞ����!,T����������Z'���n{�+; ��,Y��A38r�'����U,�#i'_�iB�g�iG��\����q�G��#
��k"��;��s�>W "�����!��y�L�2P�y�{Oǧw��w�h�6���M��݉�2}�!�xM]��V*QXY.�+�<�\����*����%�0�-ȯv�xgvkM�\˳Yʠ�U7�c�09{g�lq����Zt���n1��I�y�����ԑQ{~Q���F�1��Iȩq���Z`W�[��X�?)9W5�����	N?�G�1IJ�Ô"�T]��%2��۾��Z}���P&P�����m ��YH�쀿���o�8�ù�L�����0��n髧�{.�4vk�2[��rf��K�m�G��éU��z� �^�����+�y;��J����k��^�}Lm����(���|�vZ�cul\~����V'���;�����i�㰆6������8�R�4��v�D�5�·�a����$���v��Wa�����b�Ӱ��!���	�m���s����Ւk\���>����Q\.�O��8�f��_�Jy�E�%����N��/���Y.�3w�Rp�1�^�z�Pz��s�)����Q3 �mdc�$��X�o��:��23`��m�e�8�m�Ԙ�/UܕM � d`�u'leܛ�b#�P��r�8w��<Kp�$Eu@�	'��/��T��	���%%'G�Nxȹ�0}����9�ta!>q�oХ�����/�w��i��LNW�ŹDϽ�϶>�=GIf��-��߷�	�V��R��fx�UmyW��a��0B�)����û��q���=���c�=�342�'�X
����I���4��t��<�^��m��1�Gwf�nN{P��-�%����;� ]�X�Lѥ��j��Hh�ʟK%
?ѕ�ۋ�:��t0}��VY�2[8�=>`�P+�I���ʫbķ�!�)Ik�qd{j�����+���]���I�ҫv9m���ۙ ����w��I ����i[�ۤk�Ui=��.z��������	�NE�C����/��H��k�z�]����e�U6 �_,�w�(��s<>b���3��p+ft$	̬��W�ё�5�ʱ�s�f�'�@�,�"���h#� 4��}�x��U_!��Lyܣm���.�E΂a�u�m�����X�L<aɶ?/|,&���r����|i�]8&�Cf��P��|kD� w��P;��з�σ�_<�=�.
�24�t6
 -�vţ\3���t�+����E�c��賀G��DDC���.�Ou�a�u?��� ��C����;?��<[�8:��@��v\-i|08ڀf���8����V�a�{M�C��!�1�F+��:՝�����1��\F���*Ms?�'� ����������=�/'pY� j29�>�ym��N����\q��%��I�iz9<;DO�*5�#TI<`�gs�+���g����9\+���w�g��g������$���~�5�i���b�hZ>E����J*� �G<}�
\���n`�2ˉ�>�D�C?�o��2:��W7�6)Hz�˛g��6壢��Is�-�F��F��Ee)vS��eVu~��c�[CI�d,��M�;�d=�6}ܬ�X�GZ-��o����իg]�e%hzM߇��ѹ>~�f�}�VG.��P�|�:.���hٱx��<�S�H	価�XS�6��y�/�a��w��J��c�خhq�8�#�Hȳ��^��.��$�Y�����|���)�6!t���nLː^���K֧ ��^_���k��yƯe���A�/��IV���piV������Kx���� �^�V�>��C_F�*�Dov��*�"l�e��-'���gn6����n|T�&�X.�<�<x���Gģ�!�R1 �Ѥ���xЮ�H�s�ۡ7�=�Ơ���O�,���7��0��t,�|$6C�~x^�c�Y�Rf04~%I��\%��:�`�X��<sqgN��gƣ�g���9��>H��S���y@��ܧ�c�C5�u��e��\�w|Z�L
��t�j��A]��Z�5�]+�g�����5�ڴ� � -T �}<�p�9�ˣ��R�i�U@��ך�Hq��yFum��F�׾��B?h/Q��*�rM;�a��>�)Neԯ�>�n���f�>%ʂ���\#F�{���`����^@�Hy0{ �V�u�P�A� �h��)�9�Zt���d���tE���"����+ܫDY
��??�D��Jx�W��{���������!ٙT��!&e��5���I�G59�"ݥ��/'�(?�E�+v8K���MØ=\ܙ�� �|�(��`�DX���\����dN4��%)O�29�M�9�O��ы!���-�Ͼ�o�����(0�}�G�Gz�	(Q[2����-���x'��]3Pl�mhs��t,t9��A?큷�P$��CE��|�B��]�|wj*
[$�.�%��qnC
����T`�E r���gv�T�V���}���V�Ce�\�� ��{w� ��1/�\P��Z���I�����"����+ޥ���K��į��r��LR�E�=��݅y۔o4��,���#�ʏ&��q)Ր��ҵP��x���֝�t�����t�O2��X4�H�o��u���X)� � �lRw:!�q\+�$���f�8��h�jb������x��J"t$�q�	�:���oH�z�5��Dci�&7PL��'텃��������ȃÈ]��濯^�lSl��6c���tt�`��#�ܹS�3�3͢��C��Y�\o�y�Pz�x͜>#��e[ޤWG8���y���B0�|�$iy��w �wR�2<MC2��
�)D�����0:nf޺Y��a��G|�oY끟�T�l���j-�6;���뒧�.�|R�l�Q�����-s�L��t�m��Өբ��t:E�0�c�K˫��2%]UK�>����[[�J����{�$�y� �}� ����/.I_dl��\D�G-�Eg�2��c+�1�>�ϯN��3qTx���Уs���i$u?B�R�QQ���x9m@�Q�� ;�b��$#�Ą���M8<|��������c�bk+����s�ev~���ه"��S�v���*��`&�if@��;->0�9���gܢ�_$]5cbP!�J7�_'d0�c����z
l*�EU �k?���*AM�툊XG���S`��9�Ej3�`U���
${඀����IŲ �2�p��dC���������iD�!P8�d �h|2�w�5��dgd+};9ȭl�=�{�����p����i��u��.��~\�*�zJy��3��ё�9�p� ����'�M�E���}�a3�&�����`9�g�#o���|��6���1G�3e�����mb��^ǈ�Q�9�I�ؿ�f�됊�a��)<x_�#^�1:�4@�j�$s�[k�ٟ=�cK�Au��"R��t���Q�=�.J�mk�aml*����:��,�9�	e،ڰx����6�z��ʢ��[�ę���2o�|��9U���/�cy��]����"���ӧ�� �eL��J��rMs���j��-�1u�y��;��M���5�#4^��C�"lILk�*Z�0.L��f�S��� �C�����Wz0���A��2/+�R@��\tC@�Z!��w4�M���uk���6Wl��eO��0�\�2�� D(:7*nb��t3H���Ƌk" ����YA���`_�P�>`��|�:r�<A��qRF��(V�V��r*���g�,e�;��U���10kT�g�-_�	�/ql`	���`���l�� ��'Ǆ��/�|�D��f{�Wi��A���+~��e�h�&P˜�K"/(�U���vH]�6b����i���wٮ���>g�1������g�z�g�LDg,��Kz7�bW`�\t+4��,�)2@F6���mB��!R�h9y3��R���
�z��;�Z�<(�I7(+;߁/��~�D���\��KY'���������\��Dk��Z{B���=��7o�fd#�2�	*S:J�`MB+����-}~.�ֶ|pD_�_Ut�����Y��P���}�ί�P=�DAfkx�V	l�CZ�eRa��<��	��Xw��F��[�F*j�~|ۊ͓�#�jc�m����C�S��oʍ����I���m�>�-C�;����+����]���<cڈZ�^�f��ˊ`��1�eU	����̔|M��O�k�RՐ+k?�㗨��� ����ڀ�	e�W�e�i_�s߳|_�\P����[ͺ�pr��)=IO�ޗ���nyy=I�dB��&_��ٮ\N�g0�S�M �޲~ ��x7�U�/ʇǖ'\`U$��r�]<��`D�}���g!R45�x����3�����8�	��pɗ��Jv�� ���MB��i(hI�V�Q�(��_���wX�ccl=�����y$xnAV��E��쵊 ��y.4~��h�jQ6�i�
�x��K�/g'�.�����0�cv��d�jjg)M�|�� ߱#0*,9�f2���dr�0r�a{��Ƨ��l0h�\
��I�ƛQ>DU �r\G�yQ+��PW�� ��}C/�|���"+x�Lk����pS�[��fb��
����v�K�ꘛ�8y�wE�	t�-��~ԉ����$���%��̖���M�F4`��B���<�xe3��5j�d�����b���r̩:�L�a��o�;I~�M}O�8���=i�W�.�Х��a�-������Bk|�A�J��\���r�\�{�J[J��k�S5`��欯�q��¾M���,�l�����˥`uY�'��=�Kbq:�+��!sD1qT侟��*����� }Ea��f��En���Wȭ��ucE�5�+r�������1	Cu��fԱ@5au.��@��F*ONͬ�Lu��ٓ<��r~d����Ïr~�`0I��
�^>V��	�����9��a8������5Dr�ۏC�#�ހ�G6}�yP {(@�mY}h�{���k�o�$ӽ����d��is�?vd'Cѷ^���vP��/(��jÙ�I+�T��yJ& p���N�	��R�I��N�|[p��p�R6w�����Y����Ǫ)w�ΆE3�4B�Ѫ�0�s?;]R+�pS�&GS��
I�𐧢f�\m�kGlT�_����r�Z[0�"�8�\*�=�Q(T��Ė�Z�~���M��GDj(���{Y_��s=}G���|w���BA���\���W �WHi�2W�[ڝ���h#�C�}/��<��EtK��ظ�}Vv1�š�B���,tC7Z^�ϨJ~�� �I֌H�t�L�k����gW��XK�3��nB ��M�j�B�'�k�F�穈"�3hJ/��%EƟ�&T!=�����~�;f�!��?����ؓ� L�r3�^��~ز� ��"�r8���}=_����xHÔ"Em�`���Zw[pq�R����D�dɹ8 *�����I�*�V��R�__^��opˠ�JgMt�3��[��3=�:�+�ŵ���)���߲$�XY8��9agf����j�ԫn�����/B�󛾇}sRu�}C�iŃ�5�����^�� =S��4zV��<��_��~r�BEYega���3��~W�Ǚ,`J"ѯ�=�쯯f��!��&�hGt2����2]�������F	D�0�����6Sǡ` �1 	�;!�7���rPa�݄7E���tͣ��	7�`��%�b@���M9yJ��pa'�]Ē���Ɓ��@-~���jV"�'P�c����4r��}4�#.o�{��9L��!�q�N�)	b��P��l"�������'�<�v����K ����&�:�^)�U��⯺��8�Fy���k$� χ{?ķ	9vn��[�����Big'V���BɸRu��`�9�p���ͪ�'g�7:�r��y��C����c@������]���Km
`��; ����
*:�7�!��)���s�i'���@�!R��i�·Zﱟ"�q��������ȡ��ᚓ��D{>#��9q�~��g�U�c���!���v��_����8&�I�Yɕ��'bx�'(\u_z-H�WX�I�J��|}~��F�[���@�U�up�X��[R$����T�Q�� ��u��(̀wU�����֑UQ�G�vj([gF�_ٛ�+:YE%s��g˂n�F*�5����,J7\�U�65c�i��m���&C�K��5�w n�������J]��Q�^�x�sxIk����;�
��	kF��|I1�_:�^rh[�$�-� �sʚ���z&�m��C����-OM�|�v�D�d� T57k+N1<�~y�����5#V��̮Qm�[�j�3
���5Xa���;
��⥪���Kt����*�싴�0u�݈W��^T���^YM�f�S�鷐�Bj�o~yK-�5	���݂��|d�m?�
|Ƽ_&����c���4�L��"�Z��S
0l��n�U�R���a��Z��!�@BZd��B�e"I��'�˂�ߣ�[%/)�������qw9��XC&*GQavf���K  �=L� !?*�Q��6Ym� l>-���<l.�E9$���k��
��o��e�+w��A�j<�����5;�#7�vQ��b�`�#+O�p9����z<�y����c	겒�n������Gݳ!�a��a*�9�l|���I; �������=�Ʀ��%КI;�
	��)I߆��p�H��	pҖ�mxHp!3I�k�TxQ\`�I7|Ϲ`�rpy��"��P>z�d��H�6�gW����<������|�� ������釨"b�]H����g:��Ը��ǣ�.5�v	�1ϭ{V������φJ�O�c��CL�R\f1l�߻��ܕM����?c�|0����"�o;��}#�/����}	߿f.OlI��	�P^�}�|E�*�X�����7�l/|M+�v&:�ֆ�"*������}
�H�7����3o���ȥ�����X|�פȡŨ�\	�ґ������˖�`�m��B�!
{� ��j���dG�M\�2AĎ�&�dYu��a.m ��֚L��9lc�����6��PW<3�\���<mr��Kjk��Q)�;*��f�:��$��k,P]�1���^�	��0c�SU넮���`�"J1�$���<���ya�����[j��F\��|P��Ⱥ�v�;sVx,��c>V	֔�!�.�f���t�<X�ِ�T�Anj	�%�k�u�$�!,U�t����	�-���V}��R�F5Q@�W�ehj�	A�t�n����w�Nq4�/�	�,s�]�i^����}�V �ܐ����4**\i�`��ΰ��Vj3��AG����9`/�c����\�4�[<�7�)��	�'��[w��%ػ�h:��L��&ǬS�z� RW7:��#��,j�!f[2}}w��;\��c����!fe�ٹuu=i�o�`9jAk�7��hT�VG�M��jݺj��3/����}�צ�}J"#�VN�y5�g�>6�1������T�2bX_�E�@r�v�`���4U�hѵ(����	���&�q��2�fQ� �`�L�4�Q���`Ƒ(�c#:�3�ud����d��"�����M���q�qMm������rm?��u�P7���H�����o�
]���#�#��h������f9W���"6���$�AnW���V�N����N�\�)[�	�bFe��B�s����˚�@�:�֙�y��{вE���̭r��N��:7���y���;/�e6�G��������]&@2�����w���dj�g���ў�?�DDP<8lӢ�����@>���0<8o4�k���[�Fc��&i�Z��a����dfEUX���]ډ�N�et31�{Yx�˿�?S#�Bj@k@}��|����`A6����J�µ���nHlk
�6�Wb�>{�^�?�
=�?�5׀����|SA]D��&z��f�Cy�\�|�NFֲ�;sC;�۞^&Mq��	�p=�A�/0W�x�׈�ΡțB+������v��P�ת�ix�ٖ^� e�A��Nw+I�+���f҈�2�W&���c�b�(�<���5Gkbl�6��$�࿪���[�2s�m���K:�Ƕ�k�p�� <���gA�f�9%�"��Ag�4l �D��R�*�}a��r��tZ�k�p��;��r�+�P�ONS"���OT�]��R3�,�o�� ٤E������jZ�ק tt���B *�^�ڰi��J*�r��=k@W�TL]��ȓ.b�$����1�)���o6d����#�iz����g��_��N����gT���[��N[F�_�^��i]j](|w�[5A������3�".b{y�P��V�y���Gɧ�-��"�s�����&��Ԫ�Ĉ��]B\.J!����+�f��h)c�Lt���f�y�=���f����:�!b���v�T�A��#�k|�K�iP��v¯�X��Sc�k�!��%�:B5X&wQ�{1�㌇׎�/jVz7�s EޓJ�v�]�!�����|�W�9�ۚᤶ�~0R�d��nXM����Ac�{��R�!����Bu����X��uP��#g>��Feӿ��`�RU+HpWX��l��Y��b�<��z�0����M_#B�҆�Zd�0d$���Z�̗<�q�}X4���� 9����ٝ�0�%A��7''����NE�_��\�!g���)��K�f��"~��6��1���!��k��z��pp�%)[�y۠[$VitF���ߥgq��ܞ8��mQ�=37ؽR,&�W��SK�4�F!q�M�О�����8;<���#wN��B!�)nR2���0,:��ɾ�Y��%��5�J��i�7���F�B��v4�i+��:��I���CqC��{%rs:�wʸ��k�6j��"7R��Qw�2�n��kۅ����|+��v+5��������,��p�qЈ�S���G)�>��#Q���1�B���+ȃ�v��y��ab�<�u����k`e1�8���i��� �r1�Pk������L��(F�@{��N��^ϻ�Ƅ��JQYy�����X:�6vڭv�M����0O �(�w}s͋�l��#��C&�����ؙx���R:�.�s�[2B{�g�zH���}2�����w9� f�G��B	<�!�d���5��e}#=�B�nw���p�6ݙ]g��C����ua��.�e�W�H��M Ub�5�F�2\ԲD��hQ��������L3�uR_��w���`P���<��#ئ1�0��zF�l��^8�0SӶ:Y
x�=�*�<�0t���_q:��H����<��h�n�ǜn�?m��J�p��Hp�2�wr�`Ő�΀�5[�����Pg:ؤ������O{pe7�+GH�>��ٻ�׻��	�h �s"���k(K���;����h2���y�gL�d�>B鷶>E�MH�,a����J�*�A�?C�cC�8Iؤ-�ն�R:f٣s8�����w|��"a� 48�#*���ټE)>�'��{�.��#c[�
*�j���Nz'J����?�GI�7�Wf�JX�ж�><|��4a�o?�ܼ�d2i��[z�<0�p +ޣ�.�c����w�t�D�0�0Pg�W�L�:��s}�S�6x��Զ�&⻏Pd�śN��i��b؇��ϔ�b�&��7�z~~黺��{�a�7T�7�p��U�feHG/.v��i�Ǡ�Y�T�Wx8.�O�%�_֗��F~�u�����NT?ǌ?,�X�؟�?dH�&�G�
��Wks���TB�h/,Ø��	�ʙye��#l�.@c�稛O�j�|h���4�7<j\���G��U�x�bG�q|�Y�&�sWN�\�r�rP��R�S�&��ڝ�u�%|)z�YJi?.�����R�NC?�L$�k��$��f�/�3dD-.�΋�9J�B�S� /�:�%�<.�����sp�t���)�KE$�xKaSkԔ���Rz`�p�U�)��(t�&��(��[跍��-��g)��翘�kWK�c�:\M��Ys��UV 
���x�����@+�u�R��
��WD�`���xf>-�=~\��-eC�$��Ҋ�[�ޛW����S��v�%Щρ��I����sy�nϠR���JtshUnk�t7�L�i����g��l$�A��x��y�R�K�\��Lο�A�GCM�bm�?/+�]�᥉�����;���I�<�M$�.k�i,��i�6�VX�!*�·X>6S��/�B����fu6Ά@*`V��u4gϛ�^� 6�uk�c>+ +�X��f�}�M��H3�xԼ��L��It���OU��v�Tk�����T/E�w��������E��p�~���U�&�C�a4JAbԽT\��d3s�Nd�O���mS���[��7���Y%�c���{��Iz�/��{|qS���A��Ԯ�ph�&h�䭬D��|�6u2����@,K.H�*��T?P��������g�A>�yӌ�)Q]9�v�#����ސ�fLt]+��k��C���L$��{�>� �!�kKl��KR/,W.�8/X&�mQ�e��p��ˢߔL�\~%�K�d�)C�5@��A�R4M��KX_�����V9�M� �� �eP�&/��P�V���c���֫�l#�{77t�Mr�;;Bp�t~��1�@v�7��Zծ%�PPxp��;���6�8y1���G+�C�-���aMPyT����	��Ҿ���A��z���[̾PY^�I~9-3�Z��U��˧̤�$}�/�d���d��֔�d�T�Rb)�[w���l���cώ\a$�>Z��F4s|�a����!�x�:s�F���N��l�mie��_�n�P�o�q�n�L��&�Q/~z7\g�F[6�������f������ث�V^f����\L4 7'��	4wS��a*T�6:�c��cc��{j��R����k���s@�Z��a���R�ܰ���"�.Oi�B�y��;�b1�'�#(��`+%���i�:�~+9gB|	xp���.�,q.FÓt�f��_���~Hi�m���8�e��$��%���T�e��z�����-����Lu��.��Kd{Ag/uA���PQ��?�����! ^��d��(��Ǖt���Nə�'�F�i�!���_<��#N�E'��J��m��2�tF07?O���|�_�p� ��g��-��S>�~��~Ԟ�l�`��H�\�W��2�D3i-�X�&jԺ���	�S�����1ұH������XL���i A<&�o8�����rYK�>v�5
�A��&���4����� �#��D �eBF�t��+=ɖA&.��%fs�ؕך��W���,��k��L��/bÊrQ褷��&��],�n�:�ӝG/o��<B�����*J	]��Yά�E�C\��;�ȣu-�T�w�9�̇��>uQ�oo���d{�.nG�vʆ��}c��
����yb6�z�1��Z�|~��A�R�."N�qk �A�CS]E��d�=�Nq��Uv��J3?�t�!��^���a�R�����������p���t�O!(�vh�_m^y���Ȥm,9>q�/�\u�o�꾟UѮX`sz�*�� L"d�D5��%������3�կ:4� B�h{�|�#"E�����6��$a7��lv7+���4�����p����0�>Z(�7�O�q@���V��l�Rd�ʟ���Rx������_��&���E��qcH��!���ց`1� ��6G��(T!���t߇��>R�au��)b�	�}v��yW����L�9|�>cp��;G=�	���0��p�A�I��p���6�����_��1�<�q�ok���M�]�_k/$u�HC"��<a?jg���_D�W�S(5*�t<�F%梨m����qH�_eٰ��D����ش#�z�]��x��o�?��0���kM�Ah��~�ۣh �7�t���i}���Ɗ'jq�ZDY�z�#�e�ŝ���A��m.�~9���|�m���D�iq�[�U�8-	sZ�ip��3Eޅ���+�cNe����v�ގ� �q��EG�F�W��)���F-�P�� �Y�bx���|�h�)jl��S/2��Q���hS���2����3���d�0���.��C�+��t�������קlP��K�j��_,(c��|�ދP�\#=(�m��q4]��#ue>��qڟ����bN:�I�GNi�@4��B$ݹ�3t���
�������ݙ<rwOB�@��M0�5�2���4��`�C�}Nt/sAU�(J��w˶g�d�'-6�X����Z��R¸Xȣ�텼�K�y��!�M���'|Rs�S
��p9�2ĬE�m�"J��ohj���&֥ќL��*���f@FY1\Tr��gN�
D�{q-�qN�`��xr���1�^��iE�}�|� �H;��v�Y�����i�WJ�7$�c��'�k�Y�Ց�]I�KJ�����J~�LH��������-�-� ^��x��yߏO�����s���π�	gcD?��}^kC��	�A`(p\^��?"�dZcm�p/���4�)�&!�=f��#bd�����:0w���y0�����W�9� �%�DPOْ���On�D�� j�>��cj�Dg��m�c�=�� �D

'�$�~�}�f !�y�:�w�$���N�U�F��wB��а��J�#��w��FB��@�o�f�W��c̦�"r�EY2�I��fa���[�C��-�!'�Q�1"ܾ��4�ϑˠ�~�No�:�:C����X�^���.�q��G[m�0�iO��da���8:TU�����>n� Vep�!�$��B�����D�S${�Jַ܌YwNwE^�5��W��yf�N��'�:�z��`#,j;qw���vKMwM�m��|�������s�}�죌Y�k;���O]m��p�nU��YEK$\x+��ٚ)b�];��=!\������+Пg�&|��w�N�M�+6P�
��.��= >�!��)- '�}ǎ:��]tu�u�yA��
#�}�0<��Cd|x@�o�\+���J���̺�>a��زΥ�&G_K/�휦t�?6&����V��ԬJp��cu���$��G<˲4�E#���@N��[rY���*s���Ӊ�iF���L�J�-���n͐Րٻ�;��v	W�
io5+��KSx�a_wZ`M���lB�9�,�b��=�,���ʆ�(Rr�G�k=�5w��D���Q�9W�eZ�x	�v�e
�3��xl�^1��nC=�/Dj�GP�����`s����F$İ�����Ǝ�h3�5���6m��e�������Hr*Ct�"���*���J��x՗E;���gݕ�ÿ��O�#�������!A�&1�Q�c��ۆ����5l[�zO��z���u��X��oaM��"���j"������k]�[!-�F>sFfx;�<�����l{�֐�׶�N�C<X�I	�GA��}5q��8.?���a'���;�6P�,�I�8E�-�!�Ʃ#Ӹ������I�k�w��������B]F��W�����Ua[M�[��n��8-<�1-T��[�od���M�9�J�&��Ul7�#��$K�>$�1���ϻ��Xqp���l�Q�7��r�� y��*ߏQ�3>\��Ha$�r�Q�{�����pٞ�d��l�w�Y� ���W�荼j}���}	�	V|���\~0RJ�A��#��gY�����Ny\;X�B��W��q�)��e���Ok.X���s�iO�	�q��H%�e�#ّ��L��`�xeh�;���6�x\�6��wv������s`݁ۄ�x/�����@G�ӽ�*��ˢI7/����T��@�������O���^�&������������9a�?��~nG��/�ޡ��R+EZ:u�Qq'/�3�`�٠�U�@���>tiXpθx�����dPK��9��MGҮ4�����?+|��sL���Κ-�^��I
�p�H;��EVF+D�h��s���L���3{RFrC����k&��1��Z(bȚ']�P$��#ZN7��|�{�����e��ħ��I�}/�l-O��o���>%f���tζ�YG|�]�ſ)�H �������c��.�Y옼��)�s�����O<§]ݍ��(�A��A,8����%Y�5Y� p��_��5&u����7Q3
�(b�e�(f���e�@��Z"���24�FlU�y�ď�}�Q_�SO�CB�[��+K�GO����(�љ5;���/�-�种�e�F&�����"�|@`����CijИQV��"���{�w8��gҴP�\�'��4��3ͺJ���ǟ�QY�4͇VxPiï���A86�Ò|`=��t�WUb	1=��J����C������A9]��3q�P�����{�_V����0��(E�BD��.|V�7*:�Vn�7���P�[��69"��p�vFY�W�)�.��EԳ�f�b?�6���?_�x��-v��{e�++��Z�j�a� h6S����@���.�!�=o�C V�<j֞��RLݝ���?H~x�T��@<6ι>�:jC��u�;*�������p�]����6m�PO�3�H�+��Q����@�j�FH^�H�3Iᛄ���W'6�.'m��8��@��f����a��~�toj?)�| �o�I�F��/ֹ��9��<�Ɵ��À\Ӌ��K����vVk�6�ye�x��g6��{�$�z��,5w����3�w7���I?
A��� �o��¡���[JmM���Ogx �9d�"�dB�tuǦmEՉzغ�I��G�Ry*��*���lܧ��z�^w� ���5��������@�L4�i>��uBbO�c�N�Y�1֥S�Kh�xW��T!�M��Zf��V!�:�?��m���wgQi{	챁��MN�yY;62�E��hAg�EU��U}�~���$�7!�f��{����M�����߮�ݱ�����Edi�����ȧ�b�V��٠���������GSY1Cl��C�q��¶=ưd�ӎ�+��Pfܾ]�nl�to\Q��Cn(w{J�b�t!�k�Q���m�%Lh��|QB�B`N6�N��.5`��B+|Z3J'jJM	�'8$#��<+��$%�
E�
�i'N�HP����wޢ@�L�U���>/�E9��	6�0��P%��6o/s3��.�?�h���e�%����u�<7����$yȡTr�+��"��<�n,�h4�eM�u����?��T3������&�N����t�h�L�d(��=���=�\�o,��w��RNܱ������������j|�C���(L���~����p*����d�??��9PT����ƳlN*N�����A� �keU�?�e	$k:ץ��M�I�
n[�@2~-W�&�07��������}ݸ5���|���%��L5V��Ť�A���O�A���v���E��Q������pGs�0���=V��Q�gm��~0�t�_��Ò�-��3�HdaA8\6 �o=�N����Α��������++�&|NY\o�;�B\��/t��%��vd�^�h�����y!�(]aWWA\��$H!huMN�B�%*WM�M���쒦���ԟf���X9��7�Pp����T�c�0���e��.�u��1��>;��}=�[�-z񗽂�Ϩ+�e�G��(�Zx���N��ܽ(ǉU�C�g�,��E��Y�Cg".�=x�؅�Ҥ�&�U��f���D��M|�N���F+ i�{c̟�VUz`s[�^R�Pߣ�T��J%�׃�'4�IpU�=�3S(V��s�����	=(���EJy�PErۘ�Ug$�㶘&�q�=��������]$��@�����g�3�'4�ʋ����
 k}taZ��q�0tu@୽�P]7q�
��X{	�O���&��c�'������j5f'�¯z���v� 9����7-e³TQh#��K-ZN(
�s�pF0��
1�&�ah��Y�L�FW5�a0�M����훜!�f�@T��N�hG�rx��d2Pm�*{ ��^�LSzV'3��_��l�-(������f���Ƞ"\��ɯH�.�;�5j,�sBA(V��z�J�4V#��^��9�����k]��9Gp���T�H����Ҿ⮢��� a�&ҍ��J���p� 0��K�{�k�)"R���)�E"@�a 2����jc<��ۜuz�֠��/J�%�>(ǉ�HD��+et dG�~����q���!|cd���S�v�Ul�]��T��u	����q�6�W3M�1�:-�v�[7ɛ0��3��W\�6&���
�tE5�z�c2`����dr�d-Rz���S�S>�q���;�������zQ�jh�S�Q�8��F�@ᵱ�[^�t��e|p77d��K�(f #u�\T#!�k��@_:hڋ!�z�;�E��A:���Kr��M��biA�Ff�<.B乚0E����Bi~<�@������ș�?��q��s(�v�C�'�5��/58�J�N޶��ƛB�Q�����VU�W.�ޗ��`2�Ж�|�KJ��$9(��J���JԄ�,^R����_�z��2�]�����J7P=}}]��W)x���OjX������o���wX�h�OB�[7b��n_�O$(Z̧�{7��U�Q>��{��å��ި[��^s�pa�By��#��P�|�.҉W�t��e
ZA~Fy��@�h��t�� l�W�8�Q��uD#��P�ci���UM5G����9$�x������^���}6R� ��hr��T�A��3������P�~s7� ߵ��+�.�5�4�C��鵤�E���	"+���䗢�3��f�<3�e�L�'(��e�ubj$Դn}L�vr��R19���
���+��B�l�V*nSL�-��&�\d��g�����(C�ĤG-'}�����}j��=r%,���߈Rt���B��O䟓�'ty�W�2��uRe�ƪ�	:h@s�̍���iqgf.6����z��k5qz%�/W������2
M�� _��s�zDo:�x�ؘV��J^�(k�h�t,	k�igz�'� ����6�����x�ڱ�G�\�(E�����ҡ�д�#���Q�
��ف��Ps���]�ps|x(�]�֝�f��E���F*FGX��E�{�`��E�S�7�L�7��h�l��u�����wΈ�˒�]�X�}�J�F/��K樢��ڜ�x"�*}	�0����o��_	�z䄦~�73I|A`���+2��q+t>�7Y$��z�枾?e��n�K^�W�eO�Kr4��u鑞QR�c���jkS!�K#���SK�a�_b ��ޒ'�����ڪ�vr�@��5��9�u0����Np��>��tJ��54`��,z�ϒ��f��~�����ؘ%uɾ%��v*K���j��^����<���us�t���v%'D#�((���U�7Z�d=hE� #QWI��wu�NM�f��w���`Z -i�3��X���l�ُ��U.�*�'�M��0$��Cۇ\�$��Գ�㡩�6O�]��&�gٴT=y4h&�զ�:��ܙ���/)�V�	.}�Iy����@�H9��w���_����@��� ����A�@Cq��z$=�e~FJ�ӯ���-Ҟ ���|B�k͔$��s���:�ζh�G�ds���M���1����7h�V��!Z��r1�q�]�����B'�Y�y�mQ᪚��"���ASd��e.YG٥�_KK����~k��D|9d���Ѽ�<����P�u�}( m�ؼ�=(���/H��U%2/))I���h� �I~�R�q���Q��A�K���� p��9��ͦ� ��l��u����
��ʫ�����4�� ����%�z��:�]�*׺!5\t48����!�}�#����6▸}3��}��Ԁ�f{�w���]���q�MgK��y�Ok2�#�]p�����4?�s ��4���THP��]�Z�{
oYd��Z}���Qbj�ie�Y���<X$��g�Q܏G4��2G��(�f�/S���3����0HS��c�n�U�w���@��.ze�qU�����$N�yhS�#�у'��9���Nr �2?n=#E��@�7lX��39����p	z>�(��fإ}�9��Σ��)���O�� 넖�t��QS�'��	/�"0���$K@h�����jه��њud�r�Q~ɠ�٪��QZ22�VY]#�	-5��4'�\NԦf�{peSv�	�l�"k����%�߈��+y,�fAx��D�Z�^�&�n7n�\>"K�6�&�㸝����h�A�FՏ�,�q��Qi���jQ�5��R���$d�i�oy����L<c��ru��z�7�篷N������?���{�d��=Y���o�����%N�è���\������q�#�n��~�s��Rw;�T��DF����3Xn�㨝�|i�DD�T*u�ׅM�#$I&5*�cjVh��>U��H&a��>�.�m�m�L5��2�sC�Kf�`��&2���J8�]�(֣��]�o���mutF�z��v*��$m�x´m�?�}z> /ި(Y+����& ��B��N�I��)G!aȘ1oI������ּ���xŷ���F�yi�eGخ�?m}���%_z�Y���ӣM�RXX;�4�hcrr�%֒�;Y���Bq@���f?��0�ᑛ���`9N����(�&���~�,v-�P�-��_\�|�+]��B���^�.��'���f��ui{ƣ�	>.*�*��8�k5�{�$���j!��a��r���[Bݤ��,�~D�}�M	���mI�^�7�aEA��Е8�P��@���|=�_��V!�Q����0827(���a���@\�9�R����'�'%g�_�=�^�?�R`�йի��0��Ѵ��0�}\>�=����fB�B 	��Xv�I��l}�_��'H�0
�@��p=�Ϟ�	<��'���cc��ԳC1^j$$Ч�4��ج*�w��m�Y?��X�.�%��}3M���%�o�Y]�2�'���]�������'=H;t��>�d�N��2���&'�,c^ឥ��j�M�[� %�Y�cT��$w����*�c�1�D�g';Y�ښ.�A�	>�tv�r�,��3�-��/ohxT&�b,��������M�����9��۲4�@�W�e�xͭg��Wμƽ�Q�T����dR�5Gd�F���m�m�{6*d��7�6��u
"�o��:p7v|���,��L��06�G��?Mϭ�jC+�+]j�"���rb�?�u�!e|ẀwU'1"w�rCB W+;(�xAD�~5��7ݙ��l\`�d��:̒���)���(�S�'��G8_�~S�F�p�w��nߖ�(b~`�3��,���n:�YUI����$�,PqI�jI<6�&Ui߫88�UZ�A�*}4�bʘ<�.�~��I-k
ڀ�Y�a^���ߓ�?���b�-ᴪ�	��<)m�ɒhD���'t1#~� o2�i2�m��/ԎA¯<��2��R���A�R�M��V���)^VJ�^~=]��z3\z��wb�E�;,Δ*�9߬��=<�|�?qPH�������s�Nh3+������,�T�A$^Ci��O�J5�t�sF�gKuN��3=]�T��ƆLbuJ�dA���I�r�X�/�GI��]@O�)�PԈ�ׅ��R�v#a�«P�t�b�;�K@����b���Y�}���g�D����}<����V�]t��zy'dв�_�B�������-�<c��*��w�#@�hr��Ca���c��)���Ļ�͏���|�լa�NN\�>jZ�}���{�1g֓J��UeVgFN�e+*���4K�:*�h�?J���+�(��,�~��&?�$�ܕ�	���N��S6	�����A=a�9�8-�bx����Q�
�P�[R|lx�I2,�9����_�0�@2����#�T-��>e/���
;���%� "Gz��K�F�``��%������h�V��Z*I��@��5��@��g9{0Jh��<H��	�V����l|�y=���2�&z�,wU�b��ƾk;��0�&���V���'�j�D���[���Y��+�Bz��?��`S��H�9b��b��Bằra�3�1�b����ⅸ9�)�da�7�{ �g���0�(s�V�He�Gv�0�1�l��{�#�r�SZ�:�5>
�H_Ë�����S`P>�G`��$�����3#j7t�%�M�#�lq>����V̄���G����(��!�=҉��?�lQm¶sC��Uc�	��j�8�P����wr���0?�a�F��+?"�׷
�L��~���hCK
����v�@�~�
ќ����Us읎D�9^����A{(
���|Y��hYy��?D�4��Oqy�IXћ�KX ��/.r̠X���S�~#R^xU��
~�X-�zWs���zHF�z�U����K��ŕP����b���X�[�Es�u�)�muk.5��Ӓ�{��ƒ"�x�%s.��`���r���Nޭ�k����z�x��\&��o�[ij)>��u��7��b*Y(e_NN�w���_!`�r�	6�	d��eȲ^��ȓ#�Ko��d��Rn���R��0��?*��Uy�ͥ*2iÙ�ajʺI,�����hlrbs���6rA�ެ�D�{����.�j����M�A�rKmo�c!��Q�u�L=�cB�4>;�o��t/�f�j��:s��7�&l̨^C�o�'��/�vR\���6��o�*����DP���#�ӫV��^��M�������r\��	�~��|Xͣ�i�z�b��p�ڼ"�v��/�	?�
lj�1�H^n��6w��^�O�+�� !
3�^�:������o�-��5���s��?(�C��w#����5@���l�mO8=�����p^X�>�uJv�TV)�Qh��L���@6�Pr/"��҉*XM�0��<
5T��\)�AV
�K!	���\�Y��o���`ڱ&��B�X���P�#*h8��!�?��$%�&M"y�ӮZn8�v(��إ�˜��Y�����!b����:�ߠ��d��(�*߾������Ty��/
��� 8�'ْ�+*g̲p�γUZ4E%�keM���7�$�v�%�i�-�l���y_�[�˲�$����i����/����x��o�Vj�?u�}�����s�QB����� 
�k�<GK�ߙ�>T��O�a5�a3hy�����#��cr{�0��"�n� �<�A�5b(���1����}�z��Rp�f�bu�l߅�T�:C{)S126?��R���� ��1�i/W�F����M���t��7%Fm��K3tU��xz)1އZ�5�ƅ���Q	�Vg]��n9Y����D~X5u�7�BP�%qu^��>���N�VU�)����~�ԷK/��I$js�~ł�9B_�\���Xv[|=qc湼Z^�?�'��M�kF��A��ڎIUtM9��ѥVɃ�����cDF�y�ȕEʹìAd�ޤ��XA1t���5H6iнE9<��1[�G�u?'X=�"G*�Z1>7�0Oг�w�oo
��h	��M4f��Mco)d��:��c��«���>�d�:�����&�a>��H�S�ʗ�:H��Q~�1b5��ހ��D	h ��&�u�k1�>{����#�R�l)#�g�]	"��1A�|$Y�������o���J)|:�P�P5ތX�5B�{���F,q�b��r����;�xm�A��м������_����A0�O#�7C��\pT��r2��f�Q���m�Ի�m=����&���'z ��̓B�C6o��IT�^�3�f��tA��"^Qv�~�&c�V��0����35#��V���TTF��Nrn>C�������S�.M��A�k���WO���P�6bM�5lE��.0�2$�DL�-J*�u�m6ʭ�;��S_����7����Q�I���Ϯ��R�]O,�x�ۮ �6HD�'��e!gD��o2u�	�}�<� �OSOcl�ؒ1"���.,�.�^b��|D0uGy
�h�uA�gj�I��u�V�%?�#�������h��ͯ:�Ž�B�9C�Y��l���>Ř���,VۺT�����U�NH�V�3E4Zyy�������p� ��jf3A[������8_�|�UV�'�ЧCO�YƓ߽�+(r��l�q��:��ݩI�&O��N,6�|�F/DT�kۂ2ͽ�l���Z�7����§FZ��C{�S36�C��E�т���C�䊗Z������,��d`���uc�J�x/�t
��lج�
a�C��e��J�����ء�J��)G,��1�pS�T8���CQ^W���0u�'G�� ������DGJ�{�T�F�L�\ZՙY��_�Y�q��n)�gl]0�TҠ*�M�*WT)}��B��R�H)q�=�8kw'�p�mr�Fq��ʳ(�
嵚QL�e��y>2Y[�UD(��!œ\��4������<�Y��e�:�ރݷ
��f�5zđ['|����t)f ���� ٻ�ܤc	��;�I�����P�T���:&�:;Շs��9a �`WL��Q���5I�b4�xTU��oc?��t��D`�҉�A����fc���a���/m1�,�� �PN���X�~�;�Ca�3"23 ��O���WJEou��H��7`p�T~���A�@�k�����Ǻá�SF�6Z�HSXh:]�m�����0q�Qx� ԁ�1�@q�����Ҫ�.W�M�-���<$�1M@euЎ@��?,������p��m��J5~�q��,�P���?X�3���p"U����:�ǐU,�S|C�����\�#�Y#�x��ڂ_%�Y��$�+����e��0@��!�т�r\MR#U �"���E�cIH�ݲ�S����*A�1������QT�������g ��:����O�	JS�v�Ƶ̣hx��0�l��g�!�,��D��9�IWRjDR�SĮg��~�uN9���r,m����X2�跉��?���kDv�\�P̝W`+����ڦ�4��?5���^\ZYpPp�� p��c�%�g�x�{a�k�{FqI���*l�4(t���#���A��\�X�U��B�׿��?����!CJ�qM*)�Gv�Z#�au+ɮ��.���� �n�6���b�2V���7*�QS~G��`����T��#�����{p���{�z�#A0�S9�x�DF�¸d������M�w��#�z�A�$<�~�?�M��7��9Z��)�-x�k�$%�0�d�Bq,��-��_�(�lcVrr0��'H��t���	��`4��c��Z���[_���":v|-:1kNY
EK|��j�J��g"����M���(f��ǩ�Eې��O��b���Դ��l��/T~��G�	4,��Hb��H���2M�v�8���j��{g�>�:�cMLJ�ì�VU�??���� �E�^��X��w'wAJ'��U6��-A�n=@$W$�r�rnc/�g풑�����-�Dl�Yy�Na���I�+��~��ˏ��}'��D��4�W�C�������*bu�[���k�itu� ��9�c1]�x/�J[�⧋ �"#��n�_$�����-�ρ�7�#�kh���^� ��z��J�ly�^�q�s,Uk:�E�8Wz04�nų����c{=]'���3,r�pL�ǒ��2k�£l�s	fn�%�P�������C�	�IJ�Ց��:k�gc#ٿ�A����F�|�nu���U�
��;i�c"�Wh��Yb�?9��Y'J5(��Ln�	�xN����C����dI��N��^�����&
��1{[,F��S�R����0�o�x��̡�`e�����s_�(>َ��l]��U��Qx��N�a������:�ǻկ�vhL��j4�²Hj��zj���~P,����`(?�� ��T�����`���ېaY�f�|�R�DJ�5l�ܾ�dVͰ�W�W�) S�V2"�P�[=� �L���}�w��񄥤���Qz�L-(63�m�lkd���o�
�V�cRF�	�+��e���(�Ŧi��tsNb[&*��'rn���4�KT�3��;�I��h�[��Ϡ�X�F�E���BLjk�."��2W�+�^��%@[I	_�j�G!D!�/c�ܵ�=˲�Qb�$���*y��e�
|$2��M��m���`U���|G��˔�����L�c�duu�v�8���+�vm�l1F߯�^�şK�$a�a_�G���<�/к�1��Yî��i�l��q�5�z�t����'�w�Z�	q�kv��-1����24�^�x7�a�>�����GR:>D��އ�0��qNBOv ՛ody���|��Gm��ӨA�FG) �����S0B��P��9�~;z������u[�6�խ���L1����_j���η¾x,$��>�;g����B��J�G 	3�\+�;�����P�@S��t����6�~q\+}{�R�Ъjf�EP.�Ӭl7ua���fWS5�ѣ�SQ�G���U�[U�,���v�j��X�pm�~���#_�͇�1�_Vx�v��x�I �Z3=�n?(ti���{��N#�Ht����q��I���d��
� G�=��5[W�%�s�^�ό��.P��w���S�ѫ���ԯd���@�ea�EET�S��[�Ap+�Y���h;����n�Xu^��jlB/?+P{l���L0d���i�2�ܒ3�LCX�,D�Ѡ󅟜DT���RhY�}IK���x���EoZC�!Wf��y1�R�]cs	xC�7CC�ފ'&�eEZ�1Ǫ!��p��X�f�`��"k,�Z"lע��_����M�<�0�sl����i�K9�5gr��U�Gu�2?���B,�NW�h=�-�3��seZ�Z2��PgSî�P��J�0EV�F�zk!�;8��֍��g�Nf�ȯ݌Z���~��Ʋ�K3"�Ϗ��0��M�1��\����#VY�����Z�_�7Ģ���������%~�;�h�ڠ�ABo��
���p>�����bG����{ԁ��mp!�qLH��Љ��rx
�M\�dgAe�T��g��~@���������.����L��|Z�r��ܧ�d����J:�]�S�_�E��^�~���g(�7��s�@��_e��GAA���l2=��6��縘�E=�ȇj(���ҧ�I+_ C���XY圃��9�ԭ�'gP��p�q`+4�?�:$����i�q�Y���)8���7b4@?�S��2% ��熳l8�`U|d}W=�+����Ǜ�	k���͑���l���yyZl�K�0�/ "8]�hs�� �SV�SY���`��w����޾睙�/S̎���ՃO��]�atӁ��2���b�sT\yY,�ia]�l�6��[)��95��p���f���VQ�FW=�3gL)��C�$�P�s,�\��w����>�*hŵ�$�Cb��V�����#�`�>_b{eC �L�|{��rY\���|�i��P�'P.'�K�7W��Q�M�h���ރ��֢�r�`����E ��q|;��w	Ls����⚖ճ�3�
�\'<��.O_;��&�&:Jj�(��L�l�#����!�2]�G���Vh�g�_*+Է�F����ҴϠC)KK�+��Qx��淋kҖd�5��M�^����Yb#�@t��Qki�\��af�o�0�Rw~��P&��l�΃՝&����<#�d��&�Q�d����?�� k	�,gX�鑭5���V���w�Dx	*\�L����1����J�>�&Z�}��MjY< i�ƥ)�;������q��5<V.���������mskr�=�0��.��u���s�U��.ˠ�ؒM,4;�Խ��yM�������C��hc�W%ͧߎD��;!�7��}7Vͩ,c����U	��	{\8={"�d�3a�Fc�5� *m�^\&�_���Ka�~�N��1}�I�45�ρg�צ������Z�d��@nNR���>�<����HU1��e� ���ۗ<x���5o1#��TΛC%�&�!e'�|S���?�`I�6�K��/k3g(���+���~��#n���d:�7�ꎯ�������G
i$��;��y8(ݙ�CuY�a-t�BrA�6v�-�a�ȝ�n>�!�EM���U�""��6�k�d����F�e��B����E�m1,�n-nW���������v�cń�|�v@ E���AdvA�ӹ�ڦeE��k+���ki�O���[xNgء</��q�퀊uP-�^�u=>��Z*� a��\�W��bQY0_8�7<�*3,pز���s]�M��Bw�nUT��X�;�^Q1��)�Gv���M����6oC��>���`��ޮCQ�����IĿM��ϑ[������]�}�"0�-)Փ",꾚�Y�bdkP�Y�ky�ڡ��J
�FE��S������F���1*_au߼����_C�A����;���I�ݠ�c�'u6e���&����W	\�tEX	���ˆ�ѳ\GB,���X)�S?��	�����,�P�b��6�I�,i����'P�O��!�g�8H'f̐�� $�����-�׭��%�@nG�Z�hKRH���H��!w���6[�>�����X��{��>C��2�՛���X���`�V���-?���9p�,҃�])����*�P);C��
�쨋T�~r���/��P@׹0�v첼��AϘ�+]�
���*^̚��q��5І
'�3��y�t�ݾ�/��kPs8�Lӥ��K�T�
��9��c��?��ٔ�bx����h�I�T�H����3�F"�v�T%��Gۼ�$tζ
	����g��=���MP�~��E��YpN��b�K/{��B�8ԅо�l��գk*��F��9��h] |Β�[�����s��ncᔜ���/s����Av����a��>����&�l"w��$���p��w\�X���T�o-B���?ҬY��I��fF��f�Q��)�^����T~�<���ARۥ�b�5,yzS�z0�)_���gq�K_����ضk���u���`K�����֙7�1^�ζgL0�F,K.��Q��Z� 	���J�@�2��NPQЍ47��m��N���x���[V����ա���d�Z�{-[�pb���3��刐^��p2���ph�/G-a�D�6r��J-*Ag�_�g05��Y6�0�F����A�������bEQ��5�
�\^�\�$2�W�{���0U`xq�&4ȶH>��eb�FW��tR|�`�K�QV�+�c�|J̈́}���G�W$9�_ச{*�_�'1�@v_�9�%(9ոX6bKy���\4e;CBȤ85����3��`멛Ӵߛ���Mm�K!L͂��?~@A�$@��\r�Ⱇ<�~����[l�
֕���2���	zl����a�v��<��ޜ��-�8��b��8r�q�n ٱ�{Q��s,����%[u��8K�Ѐ��dPQ��}���'��C��L<4��`)�qu�'�[�&����b��(�����-QO��s ��o�ܪ�%���^A�)q��q(�����6|�
��v��C͏�I��Tk�$7,o�
�9b �Y�h�@0*�ٍ�2��h��E�V-
�o��z@i�K%�#�fh�ܨ>\!�.FG^��AN2"J����^�|g.��w����c��!���*���S�8�5�!�q!���9�J��-|BaN�@J6^]�s�&�z���GQ�еy���RD#�Ja� s�!U(�x1�����οd
��*d���Ԧ��t-xyS>�w��ʌ�$è�_^�W��Ɍ�P�?2����9�O���b:������^���ct-��^����յB��E�i���t����_�6�JdO����|i}ŵo��I������a;�O�0�<7�-�K��.�K^�(�r�ߕl�i�DJ4�t��9��*nIcۍnS���a�.��-��yw�{��S�QPD�{�����A3�r{h2T�`�46_�\X���R,�G����ڄ��)�.J��]�3]H��� v����n�,�M�Iy�)g��f���w�A2��K��r/ֵ��P$�t�	q�MVk��1����>:�h��Ө���ӳ*�����9��Լ�4��r�* K���R՝�cz%H$kr�7�ZPo����`_3~��Q��7��僵P!AP)�8�m�~bVT�c�s���",\��q�sG���eG&@\D�M�Rg~�cB�4̾��u��H-i��C>1_���y)I�����l�����kO�2�+L���PfɊݶv'� �����&��0�7�6�8b)F�B>W�k�TW�����wi��h��u}��iꕱX�X$����Tv�R�튐˫vD ���"��1�*���W��?��6��M�\?���*��B�^U�v�50�}�g9B:3�܂��#��Īt �h�I��GI�*��ڬ�2��K��yQ��*¶&�Ūͽ0~bi'{X�JG���Y�?�`LoD�n�ހ7�:{&����`���J�_�&��4�'8��ݮ���՗@��O�����h|6��b�;�Ώ��v	6�d�oM~��¢�)��޾w���j��KC��*@�\%Q_�#]�?����q0��l�L�����Yz���7"+�0 ��L��
�����&�B�k��aBkQ���6����a~yѝ���~M�� �k�#�,N�8��1@��A�F�ۈb�^E������9�<��J㥢V�9/6}2C���^)Y���:硰�U��f�磜�jc��17��(g�f�rc����<����*o�sB��xݣ���-�@���
��T�%g�$`гA�y�U�_O�#�)E:�A�ؕڪ��G�&�H� I̔B�;P,�F^�]#;�������&���֣+xǌ5N�nO�nE�����@3�:�Q���2=#8�U%��zKC�����d�i܈��&��V�7��{Ch��>�8��/;�fb�A�dv��.�feM�2��UHU@`���`�2{���ܘSu�b�1�N+b��^�˺VAU�0
u!����	�ʅL2��Ur�������R'| ��C��j**�����f�l��fvHTM"��W�}~?gkq"͑��7_$�@���5�csA���R�.ī.Xx݊J�H2�Nˑ�	Pl��wH���!�k>���3��7���5E�*���V];�g$�,I"��TU=�/L\��ӯϜe)\�{V4z-����z��[���7���_e>Δ-/�B�<蒙J�/0��>9=�5Y�g�쪳��z�L7~2WEC�|k͓����k�Y8,�ŝ~ig��FP{�*�!|M�.W��M1�����ujbu`0�&�ڲ�VT� �E�����\6�,���F��bR����.须h�_@���`�FB֜M?'b��j�����m���9%c����3L{
G~�L�����q�2p������+�
��33�8=��HnMc-7?�4'żݬ�N揜�?Ց�5���+�2�˗�/,�0��f��0y	5�g��2�9y6��hk4`�if(w�d���;���[��˳C�_)�T�kWe�Ӆ"Ĉ��m�,��2��^ �
�_�`{)\���j����zjȨ�`��U5��'�S�AA(�������{V�=��|��3�;n(�Q�O���n�m�55(�u@�vFnD��������?X�{���������괋�!Sq'4�l!��^��y��H5����4W��S������8J�i4:��*91�mu+�Rn1?r��;ӰW�^��+f�V�A�諹.<�����J��I��)oE=no��r��	�`��{ȷ����;�^D;���v�\V���xW���8$�ȳ�,5NᲒ�\����+�)f �C�6�U�����A��P�]��p� �o�U�
�C~����캎�z�n�ڀ��̵�Hx���d�gC3����Ϡ[�A�L�\O�� ��d��z��&��*;9�jM�U;&��z���
^9�KW䵝��u��o��>�O�(8b�H��z���ط�$}Qv��K�pD٥8���v��zT��)6��s�00#�.4��ݭ�Zw	�W�|�W����IZ�q��v:����l��aD��l�Nd[�D�b�pTrdNs�e7�����N,�Z����� �?id�K�e8)��?�f��W���@,˵��N��L���W�oGDZ��Rp��o�:r��ٗꕥ�%���&�&B�=��b�0�P�D��3��y�\��C <K�dA=���g��ԁJU��[氕���T@��:D���Zr��YVHߵ�;оP
��E��^��ũ�% /�h+�V�b
�3/�Fz��,�"l��B>e�SC7�
-��s�qBxl2���������B��,�=aP����K����tc��$��ٙ�z��}�Ĭ-��ϛՏ��P~D�/�V�]<*�4����s�W�J<)S-p������%�`���
q�X���O�5�B¦��q���D� �Rvn���}.|��@�־^���[Y^˨�6 ��6�(��b�ܺ�Ej�8��A�ч'}gh�&�y��wƑ ���@�1�	M�w����E���O�w9e|q��(�P�sio8��.qK��*�h��&���|���91V���8ʱ@�^�[Y����>ă~-{�S�};�y��0����1'�.�&�����^�?�%h�}��E�?`v��P��78eWD
�v��8`��w�[K��9�M=w�6?�	��o�k�q]��@���ꔐ8]�C��Kwv�ZyۥV/&s6NONu�<���4�D�Z\���{�a
z<��uG�*������vۍ�3:�I�g��U�cr8U�/�$HX��}����% �1v��S	�>�MRh�#Sk�c�F� cD:����u�T���r>1+��7������6)H��QMn��<�|v���8j����7�,��\��J��P��������?��Z����Z�k���]۳�j��՚Wc���)�e���Gw�M;�XSA�Y@���� I����3���1��Bz$���٭oJ��?f2����\$����`����>KP�G��┹��#�=U̮�[�.2;	��K��,�}þGe4�x@�o���aj��Teg�[�"��[	_���&Z��O[ b'�(H8[�V�c�O���-�kSL�:Θ֎�V:�"K�|�y3��e����B'`t8!�p�Dw�UH��}��r��1z����ES�t�H���٘�X�#v�F�r�Z1��!)iÞg�����|�5런�t�"���Z��-"z&,7� ��O}Yso�n�N>��������o�8UI^F~c��s=Z]���� �����K�)#=�h�L��XI:tB�@��[�c�R���jFi���'�xS*A�.?��S;�3�C��)�9x��<�eUb�w��ZH���I5PT1jňHִ������	�h��\�E��!k蟪Nr�h]�F<�Ťˢ�o���`�|^Zٯ��}M�M�+'ώR��CfG��Mt���������^�c�0r�e���q?
S�%� ���)~x?.��q�a EIp�J4��Ѻ�Y�Pa_���|X@֐ΚmPZ���#Ed���B�Ɵh�����QH4_��ct�ew�V�^#h7��%\���!���|��sD�S���d�p�Fl)y,�W��	��\���wKd�-�n,��4��;����)�SŘr����"�n}���ʮ�wb��}s�S���M��=��>�?)��Cm6�����3K�b��6dl
V<���ۂ����YC��8!��bV����#���!�I���h>8�"� N��`�	�� ������P'ͩ��I�`���ha���V_��:��V�)x9�-���3�L����BA�UF�LPk+dIF�&A4�9 �4˓��
��^��/�U(�_�S������:��G5"B���?/���˙=ʉ̑!�8Q��Ae�N�Y�c  "��G��0ln>0߼���vǠ�~o���M�l��������s�A\��h�	�B�m���z��V�b���(��̟�&�T��\̱��N�Y��5�>�Wuc�pK)F��c��<G]U]��Bq��b������3}:�x�/~W�O���e�u^2��#���Vn��h�Y�CP�s;G$/� �9@���������ȄY8��u���$�<�|t�aʷ��vẪ\��ŲB�O�^��RK���ي��3Ầ�������I�v��|�l�8?�ʯ��&�L�,�c�n��/w������}Xϙ�1i�&LwQ>v)'"k���qu�����F_����ZF����E�g�Hc�g��m��V� ?����Ga֐��e9��b�9�Z�������v�#�Š��ߚ�C'<+e����8�8�U����%�'�L�y�߼o�"y_���QZ�J3��6��G���� ��n䱟JX�w|��5)B.<��'�h�[4A�\R�(������R=;L̈́�D� �dO��P�j�)�D��8�����W'�\!�$R��WTvIq�.�y��&PZK��ҴI���[E90���Hg?yM��=?*K.�Cf��9��_W��#��d��UC�>㬱ȑ��	߲\\`�r�E���7WL�n�]Kt�4-���Ӱ��pXf��ݰشN��Ͷ�2��k��|o���s�[�i��|�O�w� ��8Q��܅�6��V�qє����Ħܸ�s�;$m
��-��@,yU���� ��R:"���+�!,��=�E�Q��Y�/�����si34S�:��NEm��D=#0� ?��W�A���ms��A�V��]���x�E�x򕄈 ��4x�h��Kt�Vw�TV3+��ס��)5W�����aT$߼�a ��SV�4��yYa���~Q��=Y�I��Nϋ��3U6G:V����JJ��b׏N�G�ற`D,��N����Ah�y����ʜej���X�t��q�A**��}�N�&��������2_����7�̪��؞?���Gب�����C$f]�����*�7߻U�œ�~_��ϕg_u��B�i�,4�q8�䚲��m�-���0���fv���ϑS�7_�Se	�����sE*����l�(8��yM��"Ei��C"� #�̘X85C��4��ba[� X��4^��Y�@� s7�:�O��YBծ��j쥋������"�`Hř����*�m���"����u�-���v�$CTdcp'��>��11��4k�fж��ؖ#3�W�<`��W"�#b�oI�s��7i��굡Y�
,]��i�{��x[ f�$�F�_�aD��P�h*,���݁��;-���Cs����}���<�Ğ�!�J�IkB�]C���c���F���z�o�)��
�7I��H�c��������\q�2S�?����59��ƞjk0Kуd�)�_
��b;a�[Y��>���0s� Syg˦z�:��O�I&�x��z�A�֔#s����t��n�ˏNY��C.Ep��J�^^���� ��?�w�s�ÌJT��9�n�(�+ ��2���!:�/f~�c!�繯�	 &�s¸��tu�4�)���?[���׼s�p���X|4J�$(��z�Jk\ߤ��;e���z���e _D�U�����b���(�����4�+� Btl}g�� k�=u��ݨ>�5]�e��=����[v�G�`̌vu��Ԣ��G�_i�K�*�2��L����cF������4�u���`�4?R�څ���2�fƩ{��Rp`7�]8YQ�R)��dx_҂?�� ]���Դ�p���	:Vጭy���c�/+[]57`��<X}/�����i�s���@_���k�-�A� �s��="��j4tHj�=�� �U7����Vb���޹�]�K2�>��8�Ӧ'����>�n�ϊ�r$��;�{o+z��pinڿ��N�EB��:��:P;R�ߌC�qw�=�)d���DB�A*��=�؂m!�Fv��}��V�Ȁ�w��2�[f�s������"�:p��FP|���د�n��@n-}=�ϣh���R6�����ޑ7Z~z�?���t��r����عrr۽���<3�;�gA�C���P�:�`���Jf��Z�q9.,1�P3;�Y�Y`c|�{򟛆������"��X�X1��O��
��X&��r���HQ�9����`�\�4UY��ݡ�#�uN���m��wc�@N���#?�UKZ��?U5�Eg�͗n�D��<"�V�f��K;�e;�^�?��P�O�t*�����ЋE��K�����?�2Y������M�pM�v��,huy�"n�N< ���^�n�ʦ����^?՞�Zp&p�EV.��q�|��X��s�)Be��I�1;�����'x�9���j��[����&OQ�i���~@����u�ʧ^޲�r	`��:XS�y.i~�D�D���6�����C��X�&_v��+Ԫ�>2�E%c,-�/8����+�#�9l�)�/�RďA-�O�������a��X�O����g6X~N�s��Q�Z|%nK2&Py���yZBzN⟔&��#�8�[zzt"�ǆ�Ȁ]Τ�C�V̀��U�H�1ӋP~r_~rs�0^޺:�L�7z'َ�O���J|�*�=�Q�"���Hh8�;y�W�h��`�<a����@#(�9.��7ER{
����{!hZlm��,��;���2"͊����0�X���w��d1B\���TD�p���qk.��� �����*2��dɱ8$�M�&yxz� �Vuwy��^eŔ��J3�G��!� �����)y�l����i��2�=�j�.\�OW�|��U�"����X�ՀLt�tx�)�N2���E�sw0}���%�v���ئ�S?�a������EC�E��g<�$Yw����5�f%8!�o��)�b`"<U� #:+���GlHK�B��V�Q��O���LR�c q1���M#j��t�s���S;+�ھ��0��l�%�UsXZL��o���I?O��L��3���N��<t�a�3�x4	.�,1��P#?����^�⧷�f�&o���K��8E�|�"a~Y��h���؅me���Q0��2�*is�/zZ)�c�Z��Q��LG(�l�?�;d���B�Vk(Ȉ�R�@X.��.�򝭎R�):{يǎt]��5���<ԡ�yh���F�F �B��}+QWpR�<tO��#4|S��P�����d�^�Cr�<�!�z�ڝ3�K�n��p9%E� �����>6�un�i�Um.���]%�"��YzN?��JR�}�5�C2ڀ�U�9��	Q~�e:M���ci�9f�g�F�.���n �:O�q��L6ǘ�!%�>V"V�&4R�JP3�%r'�������X.E�Ȍ8��~G�Օ�5�!	�!mV������9�*�R&�nu�C������W|D^C5c�f��ar���q�+��џ� p��XH��� ���#���پXq �=�]8���T��?ǧ�-��Ѳ��!��;ʗD�\.P
":�n6�xqr��G�[�.�B��2~H��Î�q�*�gҺ�UZ{�E����ys�(i䵀�V�_̀(�]��w��H�%:��ϥ��le�����/���|y�6��
A�6P8x�@�aZ����v�<>��p�2R�����j��n|�\��&��^>y�/��u6J5�]�Ug���<��7%1�̧$�ɞUM��M6<7򾏾�����0_-F�=�n��wu��A\����
���>��?(�zދf��:4v�vE[�@�{�p�#l�[�4v�ڊC/T0?����'��b�NI�D5��V���_r�5�9	]=n�7,���,H%�
��O3 �U�Y�'����"
:�%4�Ȕ�BD�O6�g�P���n$1G
���6�[�'�'x߬xI��D-��i�> ��4*�����z��)��'׮}�?+�[�h5o��M�w
������ڔ{���v�e�QJj��Y�Ҋ_-{Q:c:�k��E��=M�4��	TK��-KVU��{�ט�_�"
�%{L-]'� �����J�?�~}@Є�j�[�Po^�ɨZjh�-Y�����,_���]v� o���b�Dz�_}���l��A�n,w0P���w$ZoO�JވD1���k�B֒v�ą��e`:�����g�{���Y�鐀�AT.E~��;��;ee�*!�k��\�b.�H��q��fL�O��O2�Z��|7M����aXj��S��79/$^�
�G�?�����0m�0�ϟ�K��a�
#�6��"�����AMK0��D ��"�Q�2�_W6#0Z�R�af�Xt
 U�Oj��æ�]���b�.��X��L㛹�A���K;�9�z���,��4�U&@�f�(z:��G���2<�=*� ��������6Fi>���$V�	���B�A�Lhgq�s��#>��jO�g8�qg�ƙ1�p��^��+�� ��y�K�c�N4���*}�_u�7C��'��T�|��N�Q�7,�x]'u��b�#�X���9�to�Hz�������WT$#�o���?$ �B �5e�WG�(�@��c[�i����e��2��ɂ��@Ş��Td}� �bAؒ��+v3xp*��bLo�';yXtĻ���Sϗ�q��TPP�7�H%�s����I�Y�M�Ѭb
��;�V4��p��|���0���	V�ƶE����12;=�̨���il8�K��N��>7nk3�����a#@iH�¼�޴�����S��)�v��1�Gv ���IO����U�a�;ő7��~N�����i]�2z$��CU(�*�}�:�RAcP�B�e�E_$7\�A�� �w��
�g�o��n�u-~����)M����&�a\M �����wD'��s:N^;�*x���ز<�.���D�a��g�x�Z;@S%��zsq����^�a�g�_��02��wp�`�i+V A��Gz0]2`��w��`�P;(�˵��i��(:,@��1E���t�����@r�\�#7=�H�x?�(���=y�-��d�IU|1]J�s0���bqP �}� 9�����ڣ������8��V�9�E��;Lz��7��;i���V��ق2�7�.Uy*<�zT3�Y��<N�I+o�$��|<���t-�T���d�iZ7�@�+Rkm5������?�~&��\�1U@V��$���=�q�c�y?U��;(\��۽N���y��A�)�t�Z4�j�U�H���C�3I�]���\b�c��T��n��H������[lP3��̞^��?�X�4�� p�����߬+�c�F��KM�.�{a�����G���#%`Ӄ���B�K�ԡqkk����3vf!C
وi XU�@z�k�Ċ�,&��z��l7�ϢL����Z�/H���?���R�Yoex(�s ���@Nu�� l��S�F�>�j�y\�[m��
dqC��0���/�|�f�j>G̝f1٪D���.�q���S�DO� �Rq�)�b
�Ub}?0���3�ecz�M�+ �5���J�#P�+���gh,l=�j��Z+m�:{V�[TP,
�>�p����~�m����wX�r*Wϥ :�|��)T��0 �4���Nl1;
�yQu�il���M:4]�2�w������S俾>�"�������Kn�Y��]d��N;�
��[��­�ݞ�@� ����A{s��T��u6��6���no��B ���A�����"�ބv +�FR(3|���|�_�3���Z�TKf�.M�X��UD���t�r��Β��ʊ�R��Y�_|�_@��T���Cea�"�<��$T�*QHO��Zi����t(e�.��d��zߗkU����S7��{���h��<U;�Zn�M}�R���g�Z�Y����^Z�tA��|P/YZf�r�4Y��!_Q��sMݿP1H.%8��1�+��?�E�F�@��s�}&.��X����wR�^���"���/��:�뮚F��� piLAf+��X�A���D|��:1g�y�+R7��� �Yځ����&��O�������k�C�	~ZJ ��k������|�xݡOc��e(��� nc�!���W���\����]d�m�rؼ�Р�B�	����D^q�!n<;�k�8E�a�Ϋ-�جI�1{�(ë���c@�`�uZI��s �4D���b��n&�V�|�����u2Nd��٧#�N��en�H4��#8���JM��V�(�ʕ]r> �ZD���#B��t�g���P_�網�y����7�K2E�U�>�"��2�ZL��'2Έlm"�a ��M^6�-�2�m�"kZ58����fU|���q���an[�<�1�ll!�C���l3;�: 5�K����v�Yf���7����U��R�2��2���|R.r���wI�9I��	�����_�1�5��Y��!=չ��<��k*g�	{���{�2�&�N��إ���͉�F�.ȥ��>�#S�C�Yy9��2"Y��N�d�?�ӈ�'(ܮ�s�s�' �ӌ�H#��k���-�UX�0c���z�eo�sa7���~!�d��q�9>�h�!?z{qؠD�mz��h�Qeq+4������Q���n|ՒH�)���5����ҍ4<�@�b�1�{+]�%P��4u�`���G�{l��ȯ�s
�a����x�]��f�����H{�BW�3G�'�[S��-�C&��C��{7�\�̿�'��^�� ީ�����.)���ٙ�mͩ����&�r�)�L��LU�x� r�M�}�;�pRnv����?<����޺����/�����Uc�[,�2�#���ߎm��v�lq"sބ�{�s�m���I��OcB�Xs<1�aAhƣ�,�Z$uk�I/�l2�̯ih)rڲ׭vp���7�=�7f�/�⊕�1Qۤ�X���%�Fݢ��?,���<���_J87P���o	�Kh	���+ �33��cq���Օ
��P�D�(��
r]�&�e9j�9
�P�O$y�%���_�s�G�&J���VWd�[����!��z���q��KN.~���~��xqr�-o�C[���v��&J�8�--�Ӯ��L�nb��-
���hO�[�>�^dµ�((<��5��kz��k�$ُ�����p�I�!0����fZ�]�؁��D#�QN���)V��%
B��j�3��h���zҺ4��� ��
�]pzʃ���΅�|�bbF�O�]��sz��w�
$$Y�[����|�T+�xפQ������	�<�u1����^�"�w{�׏^���P�U�Dx������L�g�⎴Xh���|����6J6���0�kka���Ӛ���U+*��q޲QՁ��d��m�6Y��,D3(+:���^��k��Z���/N������1��m�'�{������a����lK�;L.�	.m=&Ż�����/F���f˯U��SG�yH�,aX�������em:�n�U��["r��RҞ4��U���x��43s������U�~L4h]����)+)���$�<6�c+��e�7�k��}#��W�P�\GY:~�J�Q�MB����<^�G63�Ā#A�c���:�kd��Z4�-��>u�X���vf�'Ώ���{�j�H�ܯ�x��h�/����*��5�<O��3������Bac%����U���x{C��꫌�z�1vWhn�ĳ�C�Ba
ɾ.u��ԤKg�UHjHJSG���H��������3P�=^EP������W��jE2"XnTXw]���'�m-J��o���wb�^�U�o���r�]�{�?����:��Y+��t?.X� ��l�e3R�ojo��6{�WE0�4MF�� &��֖�+��k/M�p�@%�=��^Yo,�.�������bP��&� �}���X����E�)6����R�%0m�ʁx��#��U}x
z���̱.%��@�+K\��z��E[O�^C�ɺ=q`/"y���k�U���$������Zδ�e�O��M�E��-�~��6��U�W��e�o^��e��ɱDKD����� ���1�����}��}��=��M`���y9o����t�p�װ���P׻1���5pl��l��S�_��;��r1M�P��%��E��կ �3�^-���hU�?���E~�z�UZ����- �UZ�Zr�� �z�s�"�ǟ����'��A��ܖ`~��z5��O�9��D��Qѕk�:Lk��֦�FhM0����񸮮2̴�o�. ^\��~�;%>ti��H!��ƛ�
S�D�59ą�jz��4�s�6��;9&�m�F+�AA5L+��	1��f�	��C$��b�"��f��y��(�0��/�	�~���-�)7p#k,�Q�������晱��������Ɇ�0s��XE&����SL�pW/]�)�T�ȮByX�+Ә�Ne��L��a8pz}5��>zc�凔�9������#Va:2"Sn���}�PN$z�{����S+0�ǥ������_j�OWa=>37<�E�N�*����c���c��1ZYn���N�X�~�^��=
jA)�z^"�{�e��U���}T<�"�T7�+ߏ�k�hDD���\$[S*�F6W&SJ��t0�l�u3Z,DHm�
��/	Q����^��. �m�J���se����-���ࢦȧAt��v7���R�͑`C��*��B�S�B�~�����i���+xV8D<n��/�j����Y�P7��~�n��m���r�UA0�,������ĶI�,!T�,`����\oѯ�(z�8�򝳹=�ΆO�G����S�	��|�I6@'��vf0vuV�C�Ɣ���F�&���@���1���f��i�ݘ@ �RH���C~AC>���r��J�DE"�z)e�Xl�0�@�j����
v.nF�l6�/�����S�X���d���h�&�ז���,$���&O�4�\��x�~�.�;[+p�)V��m�~���Ǩ��NL��b�ȶ�:$4�.�c��7����-���/�ͷ�0F��@Y�T<V+�u:`� 1����*4{��M��~�#����C�E@b�_����頫��4�蚡o�Â!xN�]�dk��6-G�r�r�dΎ���#��� `�ʮ���;�u������g�Lѕr��)5�E;��kFh�&��bV�]ȇG�>"uЬ<�*(ː�<��U��>���b��"���I����U�n�)��[ŀ�7`L]��б�A�DdQ)3�:Ҍz�0�їX?]�/5I����6_������H�q��s�h��"�׸�*

���CXs4�/�'mu�L0�G-O�o#P������;��*�W���
E��{�߯;�]5nG>�J��s����@���y��nC����f9.���$�5>^^�;�eom�PV�#��K?5��n<'r�̮�#l�f�l��U��z�!Qj�9n�&�O>^ 5Ų�:����:�n)�,07�L�D)_P�!X��V���,v�q�~+c2Y�����L�A Q[�7�w|>2S��c���X
&-�<���ө�\.�-���/{���.�w\�pWG���F�R��8�Z(�\��a�R)�Pj0��Q���*3�

���R��S��&�':M�J!oO�%;���)�ﺝ���=I�!�X�'q��P.�oS�Z�g|+@����{����Q�WT��8�a[ז�>�0�J��>vi�֟���Ui�>�j^�IJ��Gڊ��"ia�W?!��tt��P�O��K�c�㗤J|g׺�������U�ih��X�B�Rǅ�3#���j.<����~�G������������Ƥ�Z�#�3=������I�-�xD�qy�	��	#m1q�&'�m��j=JL�z�@�m�)ߓ<ko4D�h���R���Xi��ys��u�_P� �V�������΃�5���+�F���h%�K{�	�tR�
C8(��~ ���f?�s:��ʐX.˖8��,�I�+�rX肇0
J; Y���H�a�נZx���-��:�v��	U7$JE����8?����y%|��p�@��O����4e؟QЬc�d5�V�%'Cv�t�/� ���Q��/�|D�4�X��P�O�Q�gJ�GM��[�g>t:�����˿O�����iU�%tl����#U��0������?^�����t92��C���c#� �$
;9�,c��1 1ɡ�-��:��\�L(�E=��-��9 ����V��8>MoLJ�)~z���lvV;	�)d^4�gE�o�^	r���br������N0b�Ŏd��Z�M�x��(u0���)ͽ�z?��F���ZXm~���=��3����X�k�xO�����Y��HnZ��Qw�X͚a�r�4�"k��W3��"�z_�k.x�zvb��1�Ç:W��g}�r1!�)Yᅈ��m�/2�i;z��t������H���W���cj���BD��\퓇<�mX�+	�!4����w-���![PW�⼍��0x<������;��ޢn�̟u|Ң�6�_`��'�Ւ��7��4�����J?�Wspґr���$�o=�������,�*q����aA�Ŏ?!�Z���DI�H";�j"v�q����W��{��5��>0�9���W��")�������4@�/Rbn�s�!~�i�Zڶ�e`7��l/#���, ���IOIv�?Je����೺�1E;Ͽ�?�^<�;�l�WO�Q�8i��
�2��� ��a���-�=;������c�ُtD,`��!_��8�5~KB�iˋ�Z�Yu�|�
��u>��(���3���k�(��;�H0���/A�s�-�ˌ�rlW�Qd���[��i��h"T������"�[��a:X�����[���y6=��o�yJ�xO��C;8ݒ_��Q���Wm�]E
DP�+
1G��L��;5[Ξ�/R�ni����##��D�|��EK�.j�=_H�4m�5͛6MǦ<iU�W�(n���&�]��LE���Mڭy6�VH(�c*7J-�,B���P��0�[��u�V{�����MK��G�LA�}#�$7�8y��4��+�G�A���vq��{Ϛ��BV޶;���$@ӫ�΢g��O��c���ٟ��J��'�e�h���[�%d��"�E���5"�ޱtIչ�uR�
�*���%9?T��*�kg+q�����jMB�\�ߕ�0�;��1���)$�
/�)�!� �
�W��v\�:�&ZS�t&8�>z$����//G�s�\7!("��=w���T)�{cK����v��:��z��e�[�rޜtCV:�v����Ţ�n�jf������@v��hAAU&�ԟ��J�㧻 ��i�ғ�	���H4D�f2D�)"���w�P�|";t2M�z](�LՂR��_~8�����b�B��:YH��q!vdԌj:���ԝ�r4e����W�SR<�}��3�raă���>�T�0͐l
k6s�����M?iߐ��@Q����/��#��^�ǄT�M�p�׎$x��\Mͦ`1%$gxz�=�����|�'��=��{���$�V���V�I���߃�۞���*�Ua׳n 	:��|�^��A�U��é~��%�[��0���Ɇ-l;ƀ��'-�9��2�� ;�Nse�7u�z���'�߆�{�F]�e���J����������2 C>���n,�p��ǂ%(6�{~q�B!�Ҏ�RGG�y�O1o�xU&��!����\0 �(��@�J#爯�Q;%:�UN�,��4w�H .��ե�*Jܝˎ�<�'*���*5'�{�����d�zڽ��_r��V��1��2��jS���X�T���Y�j��Oev������_���7��ǤR�J�ꥳ����*�~f|yz�!֎o��؍j�R_)W	�a�O��J��g�̖��l�X�$F�qQY�2ƠO1�_��-�%��Ѥ#�+��i�y�Ww"���]|�as�Q[ ��͜��nN��I�&2Y�*�P���
�j. ��h�J�ޖ�|���BI��"�(/��r��[�.zAN/~%��$��XvN��T<�ٻld"Ϸ���2��R׽������姃��e�-;�U�#�e�Ե��]�����j6w2N�o%S�G�_�EG�_U�s�skGtL+%"m~��٩�9�%�7B�g�e}˥I7[����u2�BX�.i��fF3���lĄN�'@9��uLjo�4\���'�&7��~t�Nv3�,�D�$�:9Wf7�M��d��N�%ը$�Fi�zK��h�ȓ?�d&&XL�w��Ѯ�c$U	�1z���d��}M�ϕ�W�!Xŉ;K0��\S	���Ly)B(��ד�U@��h
^��j�R��3Y�<� G�������r|܏��h�fV�����A�Q�<��HD�>��x�M��<Ӳ��Dc*�%�&���� WZ'��h��x���������(�v�i�9���=�>&|��R)�/NJ���{I�9�� �mRi��ֶ�3�o�0�����S!9���I 5Bk�T_V-,u۩:K%��e�����95K<@���J�B���q�}lܶ7~��^�~��9�J�+����Ƌ���ly6kO��?��к���w��ŊJ�֒�D��9�( M��6�KSb��y����mg��7���M�#��哛�.��X
C���vR,�u�����>b��8��Rs[��z�`)���6���#U���K�,������1�����{�`i�;7��8���$vJZZ3�1�ƀ���r�Y�`h�Zx�Q¼�g�P�k���>��K��c�]���]`�ci:��*�A^�8�5=P�'�Xk�:������Z�pJ{�����=�ә��;�Rɱ��9K5A���g�
�R�k]���+�[�3��UĎ/���'��I��m����
����g�3��ѾAG��Wj@�Qɋ�8<9��r�( �Dg�>�:���:ή�i��&����Ād�=�ܽ[���c�n��ȱ�!%@���)�' �=�O(�hBE��|��&J�I�`�D��-�� ��>��3���Z���̹��?�R�ЛoG��[;2�_;�ƽ����{�ًh�O<�>�D@��m��A�2Ox�U�z#&6aR�6]Jۂ�}�M��_�Աj�N�Fb���U�<�)��|��K]��oL{Q� ���Ģ)Ρ���ۉ�ǵrK�e��D��x�/B|�k�� �b��Y��~S��SfN����{�z�׻C�N��[�Jxw�)�p�A�Eg�áoO--��u
�2*0$S9N��ҌO��Α{D C �`IOfQ�w'qr ��̿约�Q��>K�]S�B>9OG
�T����X�n��3�r|�f�	��?ɖ�;���}"
D}En�y��66�� >*[�RMw�f02AEyӐ�F��[\κ~S����
\T�A;G���:!�عVtY4�^�̓��<F]p�$��e�Wt����;ve�e���?oK��� 33�W�^r�ڄr�wj���i���%�x �z���iX+��b&1
�)������;l	6=�$X�r��S�k����f[���)u�Y���B��d����X�����a0�?��mN�6w��Out�% �a�1v�ȃ 0էI£WX����Ra�fg�[ia�eB8�>y���'a��3��[>
��}.���AX���K�{����t�]�ʵR{��ݟW����c7l���N�t>1Jr�'i2����&�w��e��	�<Ǯ���:�c�� $�A���?�����T��t �;N��d���	�z%�����G�ا(���W��qM'�P��\�5@g$�k`��I��W9�h胺�B ߊ������o��ߝ��
�k*dm��m�u��rM1ݧ�m�� o\N`��ߍa��&Y��V�{��r�?@d;Lw�L���"ߍK.�m�g�-Nb�B�D���C6&��\�G�\��Ta�8jl�//ҪZ�b,w�"�(y�f(��r�X����ZJ���F�JQU��t!=MaB͈�=Q�T��US`[�8h{������q&�貮��$����Z�n+e֒|�`�{�JcD�oȴ"�ʲ����S��8����CYIU��d.g؛l�NQNIq�d�0F8^W�m9�"f��1�Ėy?���>#JCʓ�dS,O����D9q����.K��k	��ڋF��Y���|"�sU N& �tbE>7�-5ڳb{2�����BK@;뽙�޼f6��S}��q���Yį?7d��:�����W�,����W�2���6)93��z�˄�i�aW���Ob�a��+h|�����i�{�n�P�?)uJY@�?Ymgק���44���p���H��J��v�Q�wS`QEV�3/�r�YTe���X��r�[vQve�l0&o"�vJ����z7$��/l��R�����G�u�'۞g~X����cIvN���ܑ�a��R�H�{ ޣKx&[X\���U����o�=!�	V/�b$���?�>OR%�Wu�-x�.�R<
i�,��U(�������"i=Z����]��G;����Dj�F�^W,�CڍB�n2Mo�`1��y���^hJ���-�r4f��_��Ɋ`��5&-r��ݣCԴ�i��3��߁�ѽ�e��",C<Z��qAHL\�c���6;��?�Rtqi�Q��1X��M�A:kZ`�6�\9�6|�`�V ��j�p[������P$��8��]��~��Z�x��в���Ntw�+��ӏ�`� ����%8�T%�xc	����@8��pR3�����q�`q������%�ɪ�	r�/�g�����x���gsp�9m�(5uټ�NY�"PaSF�;��l�f�����k���g�����=���4�I�?��<�N�� ���B��ݽ���g� �s���s'ۮ��d�!Y��_%fX�`�1����Z�ۮߒ�ʘ�"i6������6����À��/�vR�{��Z0��0I�]�����}[�#���H��(v��/`�i�I��$O�7����Sx b�QM8v1�:o=�~�f�K ��F���=Jt0!�Cñ?A��z۩��,az��i�_���vM���!�5�y�Z�QC���
��o��OQ ͪ*�%��Gy�l|[H�$o�s��kqrX,�&�!�ܹ9�\�t�r�n\�JI+}a��Gn�D����rym�����*��cZ���6�&����3T��X�\(�����AJ��X�/�VNܟ0*�r�X���: Y
xƙ'1�Q��h;�顰���?����2%Q��m�����܎OX��F���_k0_]桄� y��q���b{i�g�A0�wD��g������5.�1O�^��@�斟i�ŢP��M8B�Q�?�#&?�8��E�s�>j����lX����av4���T(� Y(�!M��zq���q�;hP!��	 p���@�z1Z�\c
h��ˆ�n�b�k_p��ǎA�k�5�V�~̬߳��'4����͝�L~�0���ɳ<���ANZ)��ҳ\=0v���hʤSr��hLY����(oc� ��N;*Y�^ӷG#�=��$����T�\�te�6��,Z���L0
�Q��������5���'JD��OO�=�a��@��� e[!kJ@�N�QuO��E����1_��S�{gK�E[����h[�a�H��P�d�U��ŜF����~B/\"�t�hn����E�t��꿈��i�N��[�<���6)�ޢ�pO/�L���^nT+Nwz=�yu.j�����G�=,�3F����4�`�>�M	p�Vsj����j/#J*�`�Հ���Fj|6#oSO���h0X6P�`䫇^��,���&�N�pj����|���$/� (b�-�9��QSk���ڲ��%q�U�檻�UB='W#��m�[;$-24½�f�*Ul��&B¤1��a71�L#3�׸��Z��}�R9���D:`��/'�u��(ո���rK��Qn����N���7%׻����l����2��I� ��~���?Idܱ��Q�j�֭���!;w���l�C�4���L*��W<z�#=%���?��8�����{N����ܬM[H0]릧CWrYR|��-��2��� �B8N�t��l�:�cƕʎ[f������m/���fĬ�:��*M��9���Z�ی�"b��V�L���g�.ھ�p�Z|s�Kd�{8�>�CS1���
 ��92J��!����
��\<���:�[�򃶜S��TAr��u?�6ay�"���vJ`6���yȲ��v
�3�B��CԳ>;�N��T7	э��]3�j���%��������T���/�2��	"Fp��2�È�(=�A�
Fn�I\�%Hu��D�$G����B����Zx�M�m� kL?r3_Q��ca�Çѯm5����M����Fy�`��w�Ls@�Ȝ#�gD'̓�Rʱ�ziw�p{x@2��iq��Z��%�zR-��RU�@� I��Q!@�s��g2�!aU.54�S��j�[�)<��Q��wP{���Yx�h=w@�?KCL�hk6 m��k�U�f}Q�p�[|Nϰ����(�%J��an%)ߠ{�nY�z�������jWd�C9y-�e�hJ0���
��T�ŞoDad7�\-V����Kd��Ǝ����qC�۾�v��u����/}�wٝ�3�g�z�,����x��[���>�<K��T��+k�w	�( ]H�YxV�����i$�v$�lF������|WW��r��v��UQ����3;�pڈ��lE=���ӌ���+
S���Κ�Ao�Nnظ�m�F�>A���H�l�к�_0=Ҙ��� ��{F�Ry�����^M.�����������_�$@*�ލ7���+x���n�(��(���W%%�O�_2ro��u�QP_��@#�b��$��~�ݐe�☋��u/����df�4 �/]�>�Ρ1 �s��KՅ�dA��`1�� wN?/r�`�K����_r�I��,�Q#^�^�4�!������}���WҲ�g��{�6{�ðB�+�B�CG�����p�U�7�Ӎ�8ؾ��q�%��Z�E�Xn��>q�Wq�>`[�)@K���j��Q?n���0����v�J��f�sN��@>�O��^��@��h�f�����b�ٵB7�)e(�f�;�:{��?{��aN�pW�����"�n���2��d M*�c��������I�"�z��FF���'��y�������gj8|��#zg~}<�_a<������D�#Ñ�9^eޫ�o�~��Q��X�H��Em�����΋�o����6�%�����xݨ �N4��4��!H�(6�v��n~�M �Uz�����%��gi&�o�~���W4��񭾹N�Jn��-9F ���3Y��F��l�E3j#qG��m�IK���[� |���2>��#�h�4]�g�	c*�9& �����s�^�q��ηc�c:�!�1'���M�:�-�(խ��k���&p�rj���>�K�k^X|�>��� �Mf�����"L��b��L1Rc����7�T��d�-D#\g���W��6"y�	��
ħ�پ�X��Iy��a�~"?�Dl7�p/3�>D;K�z��tYdgg�{xcUϟ�(.$�����rZ�Bf�T��8h�v��SCI�4j  զ9ߚ�&V�a~h�ћ� �0[1	:�ݬ�AW=� ���X�VpW?-eB��`��R�^DO�����:ư�x�G��dx��8���ܽ�ZE�������*d���F*P�ǲG���������hל�#e�Z��	.M'�4�������&D�l�G�KA�X<���$�a�Q8��[�3?`���*����4��6�7ca^~�ŔtT����-R�"�J������%�/���||Y��V$��Kb��|�_tG��a��ܾG�,b�2�a���&j2��-{t���l�u�FT&�stL��3��x��5�Şk�������.�aXk�6�"O�0}M�,Ǽ����2�>]��Y"��f�m�{d@��5Ld6N�i�e�&��n���hL�Nʱ��Z*g5���|�qQu)~+���"iP�
��B��><���2�	���=���9%7�J��Tl>�&��,~�GM,:�ogo��p����ۅ=S*:�R��֡���g&�W�Ba�4�r�A����})��-?���	�v1�P�4wpK�k�P��.�If�t���e�ϐa�� ?
�],��TP7X�J=��������zu�y孏�:���}A��\TY�tb���7���Zǻ����p)�2ź���̚*�
��C��
���r�|k�d�-��S|��6ﻍƙ���7q���ױ�[��1�>�͟�)|�QY�3q�σ3f®���a��ߕ�<�Q���5~� ��T;g~���3�o���	A���D�����ꃍӀ���O�T�<�O#<2�9H9��C���g��q��ß���i�W��m�*�3nE9x�f
�N{5J�Խ�D��/Q=�_*�7��KZ�e��4�>���z��8�����M3N�Wwc4a��'����W��p�Vd��n��ґ��×����h�_�J�}!��C>��.�=}�$p���;zH�Z.��o��2*��ΠX~H�����q�o=��[�wS����H{� M61�!W�q�Y݋L��'���qlX����)�;o~���[q�S�Zs��R�ߪ�|�)��w�pP��4'۲�C8&�pt���}��)a����^��b̈�hx_݌曔ĤC;"�8Ht�Y�c�W���I�(p,���4��5����ȷ*��M�j!/�؎�J��DdA��g���U� '%J�|�����gqS�s�R+c�Y�.ܐ��mT\��h����!� ���[YC��WY���&��4�����L������������J���&l�����6�����c_e"슱����T�o�.Z.Y��F�X�\|�Y���}�Ź����rG #�	g�����+1�g�d��Y�[+Vc�7��8ʺ��u�9W����Þl(ښ �{�<"eV��{4��c�U�����x�����<#lY�Ń`p�=$(q�t�Y��!��Yʷ�:O�ic��P6�.`i��,��S�b1���=�g������ �����x�-���×�H1�6_�Q_7춖�@it�������<�p&��*�!r�bԙ!�arN}���G�@E�`�M�5˿8�X�������X2��Bɔ&�s���zR��zMo��6�zʳb��ƫ��_���?T�	S���WR�6_/Xb�:qCYi $���-+�('qi����l�"��������V���z�$���ڝ�gQ��Ώ�G_������Nk%!Y]	m`?UG�D(��S�
}����?����=���(��cBa�w��9��tfG��#�N��u�z̀��B��!�Q[�ϧّ�[[�wh�}�w���i�v<hv >��-��<��	7���f0��R5OuBj�ۏ����$t���G	EX��&�:�@4P}��(8#m`Sݾ�����|�.x\�:W7Ft��A� tq1�0����ϥ��ʥ �'liY���*4����)�l_$&zj?�.��bH��_^X�O������l%-�pk���٥�/�\�p5���@/���	Ӂߝ�M��F��`�;
ɠ51���(��q��o$l}+��,�0�{t�^��'A��k`"3V��G>lܧ���%	\Vϛ����e�C��޻� @M��=���?mP��\%�3�ܘ�M�`��o��&-E�tz� ���ÿ��e[�_��o�e��G��i��9C�)P&�Y�,X;^W�O���� � ���y�y�QG+|A��	9�Eɥ��E�Ne.��CxU�a�QhAw����&����Գ��"p�(��(�܉�<�T�+�'�dǠ۪Ef� 8�*�T�������<��Nr)Ue/U�C���8��5݋X�ԃ�_w�kDOSFsɕ�e��V�ҧ��)� ��\9x��ʼK�.��vJc��~]|\�rM?6�y�u>~$���awDG�7�G��N�����.�)��X۝��9�px���6��4��z�_2.���C@�W�e>V������v����U���2�K�ЄPQ6�8�S_ߦ�4p�g���ӑȾɲ��s1v�P�ҫ^� <J�b_	^�Bsv@��ީ��!%˶t�|��2-�*��U�{ ���v��f2�I2��a�}���aW^bQ�Sr?�JA�'��3J�T�L؁��ʦ���㍵��Y���Ko��b�9�,S;�Q��o���K���[�ƹm�[K�<:l7i���}j�z���j�(+����:eg9_g�R:X��ezR>���H /�Z*��R���ǳ$Eh��Ȏ�Y6���#M�D[�.�>����̗�gu�1K������7�چ��scڻ����LЂ3L��������S�ɏ�?��v>�Vi�����30�P��N�D��I[`v��	�����2>�hWS�e��h��'�4R#y�֥͊���@��O�A����lpy$N�q�h;����=��$�b(�����<�{s�f���&wݾ����/��K0�5����7^(8k�=�Y�������E%dG-ޑ*�J��v�;�HD+rl�|�X/��4��}�B���*���/n}�\��>��Q�1�eH��� ����_�epOu�m2����z�֡
�
�����㙢Z��G2�-�},j����Y�����!&��J����S��@���{4ve�o���o�Y�<ƀ�[��a��h%���({fj&�2�IE��षS����!O�,��`Ic3"�]�VL_�S-\��RC���uZ]HN~�tb��@�*���,'�~vն]�U �l7��������jw�%w4�U�p���{HG���L����0�X�-���S���t�5or�+ R	1>]p��<8�������6��M��t+<����/������Cf�������I��Dl�{)N{}�w0��H�8��k��x�۳*����D�cbM���� cD�f#�-x���Š�81g�0�>c��C�y�E*���e:O�KA%��|,?� ����KeK	�U�a��$��d(]O|j4������}���Zub��P;�2ؔ�$�.P�95i�!������5�4���ekU����&԰��C=!��⟫�/(I��� � H ��Z��"�"�A	�Zw�������82H� ���
���а������D��b�S���Ok�n~��G7��ާ���\���%3{+��O~?kPo��1�~�!�/�"���J�����P)9ѫO��Ю���򂊬Q\�B��I%F��QIƸ���ׯ]Sņ�d�b�C�����5�fG�F��&	O����������9S$g��!�
e�������g���SYcZ)3�����T!�Q^e%��Ѝ��:�+TȬ!v]���q������]�\���Z4\���2db6N$��<�'S�[?-j��f��S$��8�����m���E1�~����R
�2�G����U!�r�=B
��T�<�v������yp���3/�� ��m�	�܈L
�IzaH�$���=5�s0J�8� ؿ �̰@�����Ka���-��p85/����s�1�����QLQ��4&��e�o�
��o�G�|�w�x)i�I(�/��:���m��-mʰ��w����-{ZK+W��q�r��)0�H�����!��#<���-�P�7(��k�t���<���Q(Ī<�s\X��i�j!��1ڶ��f����������Q��Nj�b#qQnvH�J�@�K�Faon@�$�D��Ր=��$����U?T�C�|nU̐4����F����8�QY���.�˷�}ׯ*;�&9�ʇ��N��}C-_Dņɣ����ޣ*Shq����D�M>�,��s廠�_0�KW^�{N�Iޖ1�k�?�b,��E��W2H�nm��t)���@���5Hv���%O�2|���FxG�4����<"���΂��+M(�����u�uXo)���x�|�N�L*Hh.j(W����)�1G������T6��>3��8`�x����8��1K�#�n�z)�� J��f�<���	vI�9$"Q���0�9��z�~?.�5	KQ�<-�Z��1���N{��j��I��K�m��Q���y3ST��:�	e��uV�:$�����G.�+'ك�G��s�K .�l^�z��(����h�t�\�\&�M�����Kk��\U � p~�Lj�w�=�M�n�C��a�/6�k��v;ண2�b�#C)n�#�.hDK n�������^bB������aj�o�D�<M���_w�^v,/՞B��z�9���B�[��w�\d��h=�M<|j���x���e�@q��V�>��J��L`Oa�����]�l3ƶD��\E{5�D�^i���8c�A�8�@�ʪ9SJѦT��[�:W�p�n% �� ��3 �Et'�||Dcz���֏s`�?&9`G��p�8?"($������ɣ�?5��*�d��qy��u��"1C�j�Cl��2a�g����$��u�x�	�"�9�׸�(G9���{-�B��pn�7$���wp��j���f�;_�a}Ǿ��$:噉��yw����,ݒS�-Sz���N�l��{�9�~�$90�$��m��Q���f��7�[�Kg�|)���?��@tD2�D5�d�
��f� ���B)Id��Tm���W��z�x���_k��Y�L�P~0�I���2��N����36���:@/K(��,���N�pd:{�_�]��������j�i+&o�ب�ZV���cYw�2���=+�HY����л���\�>�q�hu�N��+wb+!�@>A���7I��޼Z��m����{�t��s��/��$J��$w����NC�Er����(����N"�}̤=�!ϦY�F'�d2�� �Oqxo�ְl�G�/�&<G&g~a�A2�=�_�T:�	���X�h��6����DW$����A�z�k��W�.� ��V& �~�mP�ok�Y�s���/��ԁ�u&t���)*�w��'�=��u-<{����=�_�S�=X������v�u���-f�����`�N0!��#�|`z��lll7��@�<�Z߉�y^ߝ*�-%v��p̀m�[+��oN�M�݁��8�zA!p:U���c3�3ySW;G�2�El0W��x��o�#���ա'J�pi:�`�KT^��.�*�	} x�dl�-��c/4�>�l1����p�R�f;[�}!lBu@�~VL�̿���ݴPl�d�$�֜%�����?��,R����>��_@�ׇ���u�Q.��>x,J�L�[�Y�L�Uѱ����h"~��>T@Hu���j���\�)N��~�V�=���0�Ԙ�<�|_�$���9���k�uk	��d,�d�K���3�1�>���҃26�er�T����E;BK�o�g$z�%)��;jI@��E��v''�%i��:��N>����AI��	�̓���V^>�]�%Yg�hWYF�.��S4x10�W��،�7�QÀ�4\\�����3�J[��������69ʙ�������_V��/�q�f�ά;׹����3;-V�|z�E.Q&��E�����2�"v�H��@u2%�����)k]7% ��3{���P��T𣧃��T�,ǂp��j�߀�n����1h��M�_䥧�ѹ%��b]�C��PƆ�����9���/}�_�4�L���@~��t��L��(����?���q(<�*�H�Ʈw���3�n3�H����|e����I��c6`6l�O�/�t�};�MK���/O���O�:g(Dw���F-�\�X��jXO��1��)��}��ֱ�r��������x��hx"�|p�As/'Vm�[��X����?�QY�a���+TP����?�=}H�Sx�	��l��3�g)@i���[Ĝ�-0P��c�{�]t$[
�����_�[�bٚ�o�nE��~8�m���K��D�K�QC�D^����e'US�K80o��UP�7��W�^�F$�΋!(��f'��]�%�����N���i�s�w�-�3��4\��7�߬Ҕ�I��=�5_^
�-���W[p���%9��Y_1�a�}b��zWz�3K1b����B�J3L��2���Jl��[�`������Ij;T�t�K/П�ٮ���2��N��NУHT�dX�`~�2@5Hj�	���)���ڃJ�5�ڐ��[݉��H�+81��%��v�����ɝq�~�h�
�5s�Õ�Gb8��2V��pק͝��2�~�-�X	�lG6�"Y{�:�+��=a�9�[�9�oy�*1cE�m��i����k/���V��g_�S����tSG��]^%Y=o3��#o%A���X��P͉K���8�����ț�e�W����o��N� dK,G��g�wT�QٓjX�ň5q�Ϲ.ήW��R��q�#u���K�]շ(��1�(�5��2n>�~}nimu�c[��o"ByY�_#�w�����w(��{,|�{X��$��+LjV��R�ڟ���AGz(�s��W�^ה�G�DۃL"�����CQc׺����U��/�>�;q]�6� R/�q�?ؔ����͵��J��>u�+wR|����K�V�9�|g=Q:ʉs�YM�_�R5U$c�������I��7yն�ֆ�VD��j\�T�mw�!}D��	q�f���:�%�ɖQ���l'3���M�f�mAZe`m�E�1��UQj��d�XQ?U��6����2rG��K����Y�)l%L�.q��:�����FI�Z�^��6� v@��C�\�����ع�j�/��R�-?.ͱ8P4$���eYGF�,GK���i*s�U (����2�@�Ii	���ң�VI�?���nH3��ߑ+����F�5���~�4�-�/uo���H��+	��rZ>Y̠l��$���'� �����>���\� o9HԄW��4�U{��d~OÃ/�;I���q�w�ς"
\N���n�e��c�1v�h�˄��ޅ�cldk��SF���Sv��H>E�FJ�
7 �0'�c3��;G�W�=�:��������T��nu���J��ޝ�ݷ��ᇣ5��.(	�*�05�u�?�Ջ��)0�nZ�l����~��) KǙ/v1��|����g?= 3}�c��	�*��k�D1<�Ӗ��QB
�4p�-Hw� j�6�kGdL�|�{6��J�;��u����,��h�6l#k��9cV��ٚ��P��X�ҐbF������J/��U��[Q�f(�����ޜ_Q�m��'2K�/�z��ʂ�^�����r���S+Y9G4�D�m��l�h�[��6��-3���^�j��	�ɼO'���k��i�ԡ�e�2Fˬ I�AZ�w'����[�a=®��/k�n)�6��b̷և�����W���W~T�_�˽��:���y��)u�!�pA�@D�bo���j �<ݴa��+�t�/y|D֡��_V�F8	�d�����@��5����E=�~�,��a�iu��;��q	M�u������'�,��فL���j�S�����$���fR�G~���^D�����%�ސ֙�kp��Sh�����t
�tDH{�ΰ��{�x;T�����*`9�M�.)+�BK_.��f�!�>p(�U��J��m�fᯜ�w�.z�W6���p��ef8s+�jA�g�F.�A��+�y��,^_�@��&�����\�o�1��r�6O�����я �0�P�{4�/�{��>��}�RfO����딖Js�s#�xܥ�=�#��g~X�0 &�Jۼ�%P��T�����?,᳆�^��.���`mZb�B|sK�r��KUG|���.n��̶}��	���P;���Tt���pF2�6��'p�	v���aCP�4��KKvC?���ي3{ixAﳩ������O���.��?�B[^�Gi��Yʔ��P�ެ�Z��Ƙ�;W����	��^�����a�����7e_�Y�������?V�:'{넉�k���������� �7ce�-��m� 	)IxC��QKj��i�kp{�A��o8�%��cD�}�7��݇'�᧓��R�_����wW��r��SRL�bVe�h�����7\�-%�t�X2��t��~���Q��|���:�zV5����l��U�gK�	�+-��H�_Dm���ەd�rq1|lg�����"��F���<��,�<"�Ou*mR�M���,D�s��\�?�?�_�Ȇģn�p#�wS�v����8��|KSa�X���ߐu�zV���.q�`no�C��[�ۋ*/6�5-10ag� �-�O��w�7�������;��v8��Z���"��G���09��$�	��2ޒJ-�sYyxy ��q�l�L�_DP�q+.�:�F�Uş��O�2�ܮ��_����J�J,\X��-F�s^E'����&f���-0c��i�YQ.j�j�e0�"#����NGm]q�h�iFM�QLɞ}ҠK�n�{�CsT�ăT���������H��H怜5)`����2X�.A��m�b�����-�2�-�1#�b�7�{m�=ؠ�T��xCgXD��p^:�HzG�Q��Btg���xn��m`�hk�C���i;i�ٕ���.��S=��=:G��_a�>�
��P75̊�c�䒙���YÂ��H���A�o��ݹy4�4p֌@����@���t��t#qá������q��Ddtʁi
:FY��_� ���7͠D��V�ڄ#g������R�F���m�5t~�����co0�����p`�Pr�d���t5Ɋ��k��v�<a���W5����~�$31������E3h�Y\�D���4i���7�	&m�&��G��6����W��}`�ǱН��ư��^�:~\p��k�6�r�Ԉ���@}i���1��r7,��ܹoۦ�H�Ξ9�Cq�	8�~�v���D�ϻh�X���.���xv��C���Ð�s����o�DۿJ+��|��7��/A륰
�㲩3���T��%�����tw몫��a�(;u!R�,���л�gTg��"�Ŏ]�FY��x"{�/A���S$���-��̳��屣A�o�#�5�J~x��|{�F�i�{"�e� ъ�c(�x�}��Q�c�������7�þ�C�C���*r瀫�s͆����� 
Mm�Y�dZt�.7Z��oa�tϤMy����
e���
��Akő�c:4C��dR�7@���^��|>���R�Gf�Y�z<�7-���uԵBT.;Y4�	IJ¶x9k*IF����k�|�Ϡ����EwT�E A�e�{	e�ubj*62O��S��I�imI����@<#��8Q����C!ų@

�9�5h��
�$3>V[S,N� �+��o�&�9���eg`�Ps�2����p[w�R���� -/4cDY��.��eNn�U�q7R���BL�?�i�
���j���Jjô�;�������F~�ʩm���,�4ge�ˬ�Lr�����L�_�u�;�5��Q.Du|�z��p��
^T�"���b�D�CAc����C4�ګw��g�|2�4@3���6��?;��*���?��� }�����Ɍ.������I���5���c�Qn"��0&�'���`
j8�z�>��J�
GB� �\�kz�_����'D��棎��m��BL�0C�FO���#b��j�*��{��@���$aRĹ�Z�Θ��6��ˡ��qݕ�����M����s�u�f�)�Q�C_�1̌ۿ�u2f�<�q�T:�u�86<�b�c��0��:o:ο��g-(�`�3�(J���1�?�6��8���i���F���f����_����Vs�/��c�&�~��(�tX�	̾���o�x�:Q��0�j��"���V8�>���rP��p�=�y�g��Y�d��Z6	� N�0�E�S�zx���X>�<R�F��}���&>U��F� ���҆���crr�;��<_;�W�#G�����{�+�����65�"z(|�u%PR��ٻӾ4HԎ�OdH�,MP(?�)E����(�rg��M�+c�Le�Ԧ�L��2��64�W7�1 87ڕ�)ʊ��* ]:bl	�o��m|K�0�\��P�KJ�Z\
4a�Ϸ���l�ۮ����!4�-nJּ����_�����B��*��>�3�&�L;Ow"�lY�Z���QsO
QE���sy�̂Ow�2��}'�zt+���Y���� ����h�G�.�� �NGb�oC)89V���a�
��Ou�F��}�u_����Ro�J,#9YAsQ��jYU�� �{�$/�¥J5�0��L��[�n�*�ٴ��9����4�����W��E.,�㱾Oլ�q���}��[�5�e!+U�
�=c��N�=����A��U-a^~v�3�R��G��3�7SU�$ĭk��U\���ѝ�ATD/ɚjH1���!k"	�����'�C���άv�"T�D ����Ƥ|�o7U�\6�8P����������{+�6�
2̷�y����ǽs �����C-�I�k�=3G���(�}�.ؓ��UN΁�NUL�D!�M�#�`�c�[�C�:��V�\|� Է�ʒ�����
��&�ȷ�t��v����Ug\�HX��:;���pq�œ�^�)�'n0q��X1$�x��c�pǁ�`�L��-ޒǓ��PЎ����a���&|c��r1H|ʳ�@c�v��<�&�9��:#Gʝ��`���G�;T�C�ى4��#�����Ǝx�#*��[pՙz�3p��r�	�U�C�!^���	,�)�	�`J�<#��՛3��2 ��1�������M'��̺��ގ�oN�pS��<h�ǲ��3���#s4��-�"�A��B2���7���E(�����w�p���8�mO� u�gK��=Q���ޤHw��Z�dxO[,܄9���aA19k�p3��iI����ɧH$���#GF�ŀu�WWs11���{��J�f�l�U�xM)*�B���]��x\Z���)ܒV#��5���S�@�Ç��F�~M�h�ҥ������b�a��{�FH|0=��y��An����1hc���i|������`�&�nj�_���ȡ������.��W��=��$�h��0��6B�ٮ��}u��1o�r��o$Y�(�XSQ>N}NG,n42WVۓ�3ҟű���N�&����7��z'���	�'�Y��<�H�W��)�)�$K���k����jN�Y�@�r`s��i�F�6����k��6��@lP��A�]��}_6tŨ?ۑ��!�
���wm�G�쭚\�u�olX�D<��@�w��gqE�����pMD8V�Ï4G�g;/�D� �so=�r�1�_��g�)�`QUj��}��*x��bS��U��6B�J���c���r,��ʣE�B���+lg�D�[B@3�?B̩w%[u���^�l{'���)��
�����d����cp�zac�)ɐ��]'R�W�R�X��5C�Y��Q��$���Q���Qx۶��#Xv٪h`�H�;G`�1H��4h*�����mfj�$jꃖ���po 5!6���3.4[��2lȮ�'�9�)h��҆�T��|F��z|dF��j��R�ʍ��cW ��g�i�wC�����A���=4�척1��)*yO3�s%���%9�o+���N�j𛚜;��26VVu�
����J+銾}���f0^�{��l�� �m�~QM�4}A'@�A�:#A�2^'.?��	�h+�e3_J[L6�>/�Z7���kaD����@�|�l��ȆN�2��&�8��@,����8��!�£�H��l2��
���3T�B��˹�Y�� �D�WX���E�����6^HՓ~�aQ�ɛbW~"�qp����@?�^;��K�S�q�po&F�`C�i���4��z.�DI+��(�i��)�����p�94_
]��A��E�T�D;d��#�+y]�6����s;�6�,|�la�&yn�,�:��eJ&��F�!W�X^�_���h�-��)p�W�/ӯQ\�Q`?@�_ka �jW�t���$Q*�]H��Zt��{���Lc)�nǸ�[,�����iGpW�q�q�@:� {�lj�5��fF� 1��a6�WQZv��-���ڢ�1��\]�s�S�C�rȕ)��Й;w��$2ϻ�45��Ż�V�O���rvT�(���TϦb���q-�-He�n�(K5�l��Q<���#W��b�� �\g�mr`l��|���A�6NI'�p�P�W�:����t�����︖ͨ���>#��{i�qU�Z����c���?zg��N:}W�k�� E�ٚ�X0pJ���o~�VdT�
A�J߃�Ɋ��U��aE���r�U�Oc<�uj��o�=��-*OtU$�H`-_��2�5n8���#��Y�I���NEk�K�%���!��O��Q޲(�h�DSe�+�^�Z����-02�*�#W�C���J��'��_yO%�Q��o�]c�X�Fr����h��j���Т6��J��n�4o���a��ѓ��/o9�>�5�#����i��^�$�lX��Wk�ѯ����o��B��6;�"[�%�v�@���z�ߑV�>�uv�ͫ�o����T�H����,��m����mha
�cY_,���CG
l�J���&_w�9>��dn��iz�d[��>JEu��+�_�$'��Gӛ$M��dx�N�ԃoMQY�WzhEa�L�3Y7HOB�?�U���`|:s���F��]F�oGC����G�}F[k��7��3����>�1�
vz��ȗ�敃���
��UsO�b������˭Y��{z�uT9{��@�=O�*7�!��x2�r04�[�!�,ǋ���������8�%�Ь��1g��
.E>)|����U�L+E�(i�@Y��J�oI<���8�k��
#F]��Vq�����'�K6M��b��t�0�v�:����bHL�v�9��=��u)��!���u`{�  �@2$�&�j�n��?)N�Hލ+�v�w�UZ!|.\��4�Lt�9���� ���sK�ytϖ<�����$	�9�����މtPаZ���f� F�M>G�F�`��]R!Ǚ��g�[��"x�j\ͯ.����Bv6�Zc7MT�V��/�8��:8L���%D*;�W���P�x���<*���a�p���~V�k�"�0�,��TÉ��N�k��u
A�J�ғY4)�Y���PRD!/�Y��@�c�"�0���bUY8VW�{oq=b/��d�I��O�g��D�����U.D���T�x�d��!}��d3���6ҵ�*���;�x�w�S�&9��	 �ʡ�A8�J�X\��^SC����s21�%j m��6�*������xoӾN���v͎f9/��P+��D�|��E��}�[:�~fJ�ĵjPq��u�G8\wor���"\�{�4�V"q����z�ޘ�Fds��>�2�+�D0 "���I��Ϝk_��6�����S�UW������K����t�5�\^4@�b��j	^������H��DzA�&"�B�4��{��:=�e���B�FL������"��;ly�!)"����
�Q���|��J��Ù�+��Hh�$��t�R�±��h�m7�pW^g�rU�o��D��Dm��]�5���j!mL�>��� y	�/�P�<�OP��u7���N�ban����E�v��.WȖ�pc]�ߊ�4'&ṿ��Ͻ�/�xp1XyK�� �_�~����қZwg��¨���Ti3���y�W��d�{�I��X �E-p�M�E�gB���F���wP|�,�KƩ-y��-s��U�H?"!T~��ݛ���5Ԃ\ފ�b]Z ��&��:�2���m����zJ&K���8i_�imþ!E���qBR��,����R����	[J�No'�.�Ѱ�`^ݭ���-��gy։h��`X��Ӊ>���#��77LC�gz׫&�Áx)�5���K��me�k� %ҴgOi�j�b��L�.+���0��~��/���o��ߪRa1�
A���T/�P�~��e�*@oe��v!�@ۮ)��y�k�7��i5��|��� ��d�|kx��j�;��Q��sN`�����)[k�)�F<q��MI��/�w/��o7�)�A0����{}��p�|phV=��Gw�	��T�K?�Q����*$���	=W_�����z!X͍�5�&�z]���<H@��E��Y��h�12ae�×��/�L�`�����z-���F�S�I�%�\u���Hdux�� w���>jKBS.��3M�&zo~<D��
�*R���9���ksz��	%u����%)̦���������2{�"��(S�>�(PP��@-uI�����~��ۅ�lA^٤<��2]M���V�J�:��Z$�)��ƹ�ow"C�l&�'�����qy��ྒྷ�5����6�U'�|[a��eNv'{屝D(OW��}K��_��r���ZW0jJ��4�G�LXR#����I$I�5�B���6�b2�7��t(��*�o�x��O�>>p��ɼ!��4!�Q�$!x��X�����Y�!�Ny��c4Eoq��#������*�:��F��zA���X���0Y���vX^T;�ZGfK����,����C��Vzk�]&-����Yd%ׇ�Vk��p^��6�ˀ�⩅@�����{�N��}�D�-����Tf %�6%�`H������/��N1�� �&���g�L�>c5~��5U�u�0y�f4 j�"iզ��G�Z�
ʘ��h�NA�֐=F��</��|���`�Tr͐���w��M#	��dD���rvox�L9���/�-�((��G�!d�Y�NeA㮃�h�k#>��[&�r|+vCU�w6�y���c���G�����9�_2-�M�~ȝ �&�ef<���>Mނ�O�<�e�T�����F��,�s:��$��S��\ �n �<�$�'x�5{G��h��g�:E���b�V8�%� /���rc�36��tܭ}�&� M
Z*'�o���Q�������7´�<���yՕ0�>���P#Hƴ��"��"2��&�+�0�S�67�xAD��ю�R�ՙ���b���ݱ/���s���B�M�[h��L�u��hA3��c�ޖ�=]�y����l%.��P
��K�؜..�C�JJ<���U�[M���55��4Ԍ��1;]ƒ�m�4��$��r!��wf����.A\���Η`1�G��|�a�vT�AH5�5g.�H�r�Z��{�p˫'[z鵐�j��3u� �WmC�Q�p"�D?������(mȕZ��Ρ0��֮R����W?�9{��LVJ�y�,�V"��g��Ҍ�# їJ7o~)e񴶕u���W��K��̆��FR�_Y�@�.`w��U��1���(�{7��iE���v��fj|�	)�n:p�oc�V**0���˟�eR�"}Q��W��a!z�!�6�u�ʈ�� ܆?�9��]�
@L&�ܖ�`�(��$h�t@�\Y�B�Ѐx?��p�����V5Y�ڴ�|�ޅ���Q�a��� f����}ĝ8���'ym����T��b�F������ԕcEK��i:�Kx�/�Lv��nӶ�j2��#��|�\�ć�eκ1b�TL�Ѱ<8��L�q��>�;����f���`Hr9��ʪ�����iB=��M�+ �TZlf��[�	U����	��㆔ �p���߲�ND'��vjЈ$f�������؛��8�πc��{�mT���I�y=��Ԅ���#�_� K��)[��y�G(�U�(	���=z;~EX��`<iI�hB)��|,R�J>���q��H��2?����Ɉ��VYܳ��14'��c��=2M}��0�y徾I�
lZ{;=��UC�������K��;���%@��qy�m-���C����^�߄3ˠ6�����M�.��#%�i�z��Є��-��CogԄ�N(�E,9�Ey�ș��ԕ ELzW��!1I���s�Ö�������C�K�����W������xF���L���W��%\%>5����'��
a���4���n;x�oT���:��$.�M��WE��(V��]h��+3�+gm��'&�THC�F�(h���N!)�`H}fsY�F��B*���>�b�O��L����ne�a�"g_у�>A�-U��-e�1_���;k����U��/�~V�(v.�����}�7u�r�x2���U:���[|Xu��ǅ?��n�,����NVl�4M;ő�ܽ�Eb)n�ʨ���ߤ@[�}üGX*7ph{�l���Ou{ H���q{1o_S�A��Mu�*�����S`����.[��&�Y�v61M�_�ޯ���PN�ih���F���V��،�qQ�ڂKR�z��$H��
�?;d���Z~kv�B1�Ɯ_K���������~�����~T�'��b���-���UL r�v�+�J�5�O6
>���>=�5�����t0z��(�wn03�d��#�xu�!�=��whJ���9C� �G�@��_��@k��>G[���ђg�o����]5����X�B���zv�Yq�%��5��Kjc�X��V�Ő�D6h�b}�R,������R*<��=�Jb3�N腬:���Ut�?i�|0 b���Gg��u�G=ky��&[(���&	֞��b�/�/��5��������O�	+��a�gE~�  ��ęx{��u�-���*
[�l��4���%��<� S�>v)�������g2%C,54��+Yl��6D�aZ�{= �ZF�)ǭ�RR�m�d������ʋ/l; ����S�MI`R���6����Y��Lz�P)l�P��U,�������f�!4e��{��m����/�p�b�{tn��_��VebB\�ħV)�!�j�����B��š�a���=e���Q�m?���6�	bۨY��A�ֳ�*ܻ����8388
k�����5�O�=U���3����D�x��v;ǻ�NP.E1��I �Q&aň��vwg�'����Իu�ԢF���ƠY�77�m�-T��RH4ղ7Ce�,����I#,���x���ŧ�*׶�+�R�@.T"�,+���;"tGr���C~
�@u�P����UJ��Ac���){���u;��R2yBv@(�pǌ8r=^�fXl`�2��������B�.�D�-�O�`?��������c�~��+�E���5��X����Eo�U2!��X�¾��V����f����Y��ĝz�Š
���c�.�Hpɩ��Z�#M�hw��r]O&E{����7o2/2x��H���	�4��}9�:��PUB���BP�Kz���wocu�,��6����i)�e��fE���77��Yu�|�
�m'��r�������x�*8���Ύ�_�A{Ï�j�-�}
2tw.����!�,������~��e��@!�\���*�~}��<��t�O�]��e	���48E��m)�n�̘�\)��r�{㐟a\q�n��
�q�|�	{5�����򖮂� ���H�ވ�Ir��I1��r[ʭ�t�L�TI�;��˳�[씦a~�dTJ�|,��|�/z�W�(!�F&��3����`\
����ӡ����(�=&in�v���u�H{�cRh?�����7)$.Z����xO�@&7N�~]Qw�O�PTjN���l=a~�>ޠ݀����G�D*�"E&|"�H|�}||���t�Ht	�=m0o���2g3a�)�����Cm���۪)_���r��1�1�ϱܸ���*Up�¼>����Z�z�8d[x����d�
�jK" ��$\R,>�dv��V�\��dƃwt%X�
�h���JUF�������{Iƕ�R���������Xk�f�������
s���+�%���bE��@^ ���o���$y�g��v�,����W����U�YQz����<YX��1�_�y=��b��ak�����_�G=�Ehݽ!�E�^}oߟOW*l�]���'�Y:�bT|9����%�#�X4��|�K֔d��tDx������L� ؿ�㵮��nR���4n��Y�/g !�I��[�w��~�PB�P���,[3���͊�8	wG[� <��[��v��������Fs dd�}��O���	<Q{���Y��@o���y��٫��:��y�e�4������(�l�2.L��}{ c�SP�������F�uQS���+�mI|	,!���k�#��O�=��W��[-c�@�,�����0@n�L'�r��ng�[_��E�F������&�[Kߑp{��#dDi��*�{Ϙs@��Lg�.�H�*�[Z��xM���y���Օ�K���k�cܕ4\��)���Bco��]w|�1w}@;���h�E����D��N��A�'�Q�X� �w���r1�X�i-��9������}�m5禊�ȏ.���{m�b����Ȇ�8�㞤
C���/���5����Ov��^	mQ,�q$~��>�#YNh�@��t�uq*�]�ɯ�׽���V�a� ����ށ���-��7��񚳪�̍����?���h���`�g62������P_T���%+��f-!�dZ@��Kp��/\&H�*'V�D��F�vB�Z��������i\Pb�	��Qo
p����p��PD�F9�
P~�r:�ܩF-j<�v����w�@!Db���9�>}dQ'O�!Ƙ��޵E'(�������� n�Z')���v%���_�f0��zy��r�����Q���V����a�X����|��7K@���!te�[�Q�Z��$���M9�}�%Ŷ�J��� T�8�,��I��{PTW��.B@�=���s>��$�Qݡ&�m�]���o�Y#ă���NR�Q��(w�i�nm�\�ub2L��S�+�����Õ��(Q�ah!���-��?a.v>�
����,�u����Ժ&�dD-s�r����4�"^L���0�� pFcs~���c�(�5;&�W���f��ʌȧ�@�7Sq�6b�Q��ڧ�N�DD¢���V'�Lf`OᦦH�̒��J7:w}2�-�Oa;���*`iλ�h8zpGӈDf9�4	QRb�m��ق!����-���WWK(��M��]��'8��TU�>��E�K�b	Ҧ�:�E�~��������h������fU=��e���D�黸���Ӊ�$LK`�������zR��ݨ	Y>�q9.k�[x,>f���4[8����cx�A��%ZG9��,��ϻ�x�BL�d��xT�U�+�N�}��'7�l٥��6��������1��2:������{ۙ����m���������I��� ϰR��*g_�	��u��|BzK���p1	0"�ڗ������!�n�܎NDN�~�VH)xlv9Ei���h��6��<��>��甾���`�(�&�(ƿ@@^߼��`�>�7�*�Ȃ�������yo���l|��z��u�u�.�&�S� O�|D�$$˃_�O����e��k�9�T�qs�d�䳺�8��G����$�_���l�Ѝ�WM7��JC�W�.�wM��Tv	���˸���J��4� ��_�},2��U�܀i�>Mr���#'z\�5'���.ݥ�9��.��Q���$�<���5������i���}�Ø>w��MB�S��T��9�j� �����'�c��+�3��1�_q)�(�׶]q%o#&�	F���oT��P`���vn-k�1y#dE�(��T���5=(�;��/D�YX��=��:W���=\��tDM��'}�T����+���~C�АR���rԌ��s2�����\B[ܯ�K��c=�<5Q��D��0�/@���o��颶��_�4|2��8NV&�ay�L��p��5�V	V�/�J˔�ܳ�����8���G�흚�=6h��)8����j!�*���~k[���#���Q.9O-����Aχ����Ev�`�&G�i �sS;%�O�ȼ	(�!w3�	�2��m�����69�.{u�WI���z��Ok�pB>נ���c��:���>l�o�i��s'��q�ݦ�P�#G��We�_�%(�@T���W�v�����:��:�+������=�4�_L�[�A��v;����1�2����*Eok���&!�l�_�i�TU?�����MD�ݫ�fI :�6���OE{�� �nI�����5'��O#�u!c㴅0��9�w��%/�+*<���%V�:˶r�>d�~1)�|��Z�#%�����m���U��*���i��q�"d�`�s���G� >R���?8��Nt��b,���-)�2XX��T��X�i��:���������1�d�H�锃�	E��s�#��pM1�_�m�GxGϊ�q=���f�0���7@t��ؠ���kU'v	���@�������]2D[�
�a��w�P�]CLkYm���U�`�X'����g���fI���1+�ZkZ�M65FګW�JIH��p�.��o�|�7�c�wڃ) ���)�N7�[��u(��^7|�`�Ǹ 8���p��3:�b�LMX-��Ҩ�`��k~dC�h�O�F�9�f�_XN�/���L�D�y�?1���N���RH?TŴNU����L�_O�D��r��Ʋ��z|�I@�孋^�tO��х� �V]"�,�8	��T�?ƞ�l��$7ԁ]jz/G�&Y�4<��p��6�i�����3o�в�=$��E���5�Z�P&�&e��婹9QK�7]u�Wb��Ė���~���>���Ls���h뀑y^Iy�M���t3G��|�s
ȭIϧ�YO�U(d��^�\�%t>�,���m�Yhh6��b���c���E�̿M��򱐽<u��Z��_����!~�t�9�H����W"Y�'ޥ������/ ��o��;��eMJ`ߓ�O��!#N�RK`ċ�(	%���-�]��eMr��%˗�Z��2M�iP�ès~fX��k���RLp���̄<�bdc5�ߙK�g43�&W#��j���~Ɂ�u�R'�0
�q n^��k�`�Z>p{줐+R���|� ��b�V=I�9��3�l�Q�4#��q ��\Y9�ʻ_�^5���4Eo=v*%Y��e+x���^�)#Y)sr(Q�i�x5�UW�f��9�K��D�rvq�$���T�Ap1b�B�B��<2@���X�\�Y�X2,���2+�сN��U���3HI?a!���*L��΅������:]�-���<L��G�N
�NS���N��Z�S*�n����@3�<L�/g�.�	p�2��P�>�}_�yw7�>�|�Z�1�������2^'G��6GWR(���.z�<�Ԫ���^+2ܣ�&F��E�-RWބڶ�����PI�4���*h�}�H�3�Qޮ���w��[�l�ۛ���O��8����pE�@ [y[���h�teH�z�
�yky��!Ϟ)�ۭ�`b`���t0]d,Kai�0]����pK�)xa�+���,
�����;���<r�&�/�ӹ\�֗��y�ͬ3�eL3DU�+LN��YX�Rud���ѽ�TS�)��VӚd:� ��!��
	x��W�a)"Pl���꼀LJ_C��n�܆V^�PU�����O)Ƅ�j�ѷ렯g�H�/q��C",��x�dw#����p��5�M"�	~xn���x��o-i ��n�<��6x���k���䞣�]��������D��j�5P�h���v,a��%ىT=�,_��)p"o������5�e��hp��[q�����K^�Gwſ�%�w��E�sS�!�����>�t��5���e��,_�X� �qh��h1���$�-�
��'����~���_�w��.��-��)�Msh���-,S�kA�?��ᱞr%��]�Ӻ��Z.��j���qu�ytu� 9<�Z��kk�ދ�=�.�K��m��	���n�k� ��o�z�Y:|ke^�͹�~�=Ɩߏ����Y�cL *��ɮ�Q�/��/�6U���1I��KCZA�6�G�S��W�L�b*u}<��pó�oα�W���L��O���A�뎃�-����j�X�ؐ���C+?�H� Q�ˀ��-�BW����g��v�iS1���<�q�zԳQ����˃����B�G˂�x�����Nvk����kD3�{�������Ϯhy#�>y�hyfw�{�+����<��@�X�����r���V���ɰ1��m�q����K+��`Cv.!�Fxd�S�;cT`\66�Q���$C����p�:2����0\J�,���_^�_'v>�<��rQ��I�i�9�Ǣ��,�=op���HK�%�����n��"xϮ�j��ʬ���&fxK�y�@�f�Mm�!7�YT�������[�]ay�#	�ә9���c�s�K$h9A����S8j7�+Wo��N�"_VH&��B�M/k	om�NO%����X��	��eI���?T%����HE��.���7T1V=��g-1��a��q7|n�=��#��x�Lw�"����D�_����K2��얕��1��j:T��g ����8�k/�.���=�/�Ҳ�Mȏz��O���hmI�
��ۉ$�|�Fߓ���-�\�4�s�!G��1{�-�)?՜��b��]&�h@�d�uw�m;�6�f�O�d��vJ�&�w�����ahڛ�C��-�L�K+ ͍t���;�?ng�ܣL�𨿑���%�I�����j�;�������o��1'lЯRˀ�	��Z�#�5�����x>�7�D��KR,�ר	a�R�=$N��/ˬ�X�޸+�g��*g2}���^�<���zlJ�e-�ɹ��³>m�c�"��W7W���fYS�6��=#���}�ˀ�Y�<��}�;\�����]vϟ��~Fƣ��'d��]a��F�f�?��א�!�ȍ��r�)����kܕ�J��4���k�H��}�z�k�@��鬙�����bf��Z���eW�\r���O�K,F���%۽a�Sz���b{u4�0%AHx���HE��&Mcf�����s�,��Y��s����ؾ�϶�KIYu��C�TFHY�y�m�r�ʷU	�y��ؾ��-
��TB��m�Fؒ� F� b����� �
�����B�8�(�B�W�"��m��Gxʢ���V[뮺�_�{�W��uoT$_�,�P�����>�Uɔ��gj�7�Ǟ�gX��T�n���.,�2�-�LA2P��uY���S6�$*Ї����=Pu�6%�'h��C��B nGF�쨬��_�sW�Z!���4�����k̲��'|]��Fq���V����.E�z����~Z0����/�����qNt��/O)f<����>��.�#��#˫��ʕQ_�Wo�����Vތ� �?�q�qP�z�qQD��\���O��1�{��� ���j��n|����O����7�=`TB�Q �WA����W�}��9��RTM�ݟ�k�` �	�o9���Kv�%����Rq~�����ѣKd�?�.�f|�@R�4�v:�8�TŸdI,�5�䎋5;�2䯛�Vr�j}�Ϸ+�G���xU�ڗ�۱1S׎u�-�gj�k�z{��GϨ��4;�).P,�EKDM�̎h#�U�Pu��X�O; ��ū��[t�4&��#Ǣ��m==��=�F��0���	)����Ʌ{:��+��q�L�L�}0�@���$�:I�e%�0I�cVO��/+�le9�����t�W,X��O;ȇ��͹�㩇 �W�|��]6���)p���3� 9	���̮yJ�^^��b1�3�O��I���	����´B�z��"�3�U"*H�EB�}�T���ܹ_��s�?m�٢��A� :��=����S�j��e�b�E|�{OY0(D�S��v
z�Љ#�"M�H��X:k��V��g��B�����~%���1r?PI�C�5��lz޻�TD���<o����y�ԕ�4�YKv�R����6o.�`�/��6�	~L�&�r�6������~�{D��G�(�b)�����u,^Jxpf�hݥl�)�4?��pTz����Vy��fF,C��r.H�KԳrmN�v��j+��u$��U'*�b]X|Ҋ���:�6���.��m�SX;܇Vom�sg@�5%�!���W�0m5r�O����!�ΔӃ<S�{p;ɣ~߻�=n��U��,:A�A���Z�@��5��{�է��Ы�v����0�M+O�Έ*��NW���,�&��R�4�����ҤY������1=˭6��,}�d	��OVvĲ����Ϭ!�o��5�|��+u�b��_�UZ]�􇊥+��w�Ϫ/1y���7��r�<�)����4�^�I�����K��gY��֍��098J񥺫T�0�>��)��(�4	����A����`b_� $vٺ�8�䫓D�{k�#��K���bU��U���ly@<˗��@"���վ?"�Զ~����]�2��)�l<P���$7���g��r�Z#zj�����}��H�PP�F-��2lk�]�����_y!�god�Nq]�����g�+7v�p꼇�+�P�îY=�cЀ=k�]Z��ant��`���+!�\� 8�k�l$��t{�pq��	���"N� }�����C)98q�N��ݜ�U�������������"���z�-�\M� YR`��t�kP�M���"J �4���8�y�V��	��5�$�������z�@]	�O����vI�K�����=A���⯣�����+�;J9�s���B�L% �i	�bh��P��S,���;\Ɋ�F�p����6�3��/��[��D�6p_����	'Z�v��d�*,�uf�Z�Ӧ=D�z���^��^g�V���nt�h�3�*`b[R�\���Y��}�3vm�)���M>_��?��]����S�9�{ض��W�¤��Ya}��C�(��5Q��]3�c�N�� ;6|�������$�I^ ��_4�k+�� � x�_;���O��ȿ9C�8�