��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*�U���F�GXЯ+��;X�E	��W��T4Y�U��)�6����J�؂�D�!	���4E�5�ӂ���6n�Z�K2B.����"8�j9�T���o���,�}G� �:�xt �m%%?/ ������y�����8{7��Ų�2]�O��R�y׻��Rd���r�8���6�0q"����t[�{���W�a��g�^��dk��� �W�j�_R�i�l>gp��UG�Bg�Mk�{!����+�z��0Ҩ�^-oka%�bOH�ObP�����0��Q�@�����[R��;�������3��[�$N�c��r7�M�>pP��I��@hV����
h�8��l�]B��X>Y�C��LcΌ����""f74�R����t�<[]ܵ[ջ`���h��nO$��Co����Gm�N�!��/.�g�"���]g�|Qg+繭~�#��G<F�%/,<4��T���[�\�1%���S�4��X�r�/2�]7��'���D�YN��&��<KW�q�.�c^�I����2�l���(};����#���y�P�b�g��Bz�*,�L�0�P��@ $�]!�� /���c�d��/9�P�����K�Q�?�O'j�v�; �&I�n�p�+��6�����L�ʄiQ�rm��pY�ss<һ�a�%�4<�4��o�u�M��;^��gęT���cfD��!���V�;2�$���rc����B�v~�C����T�����Q?c��kjI�	��c�x8��:�{0�&S��x�tm�0 �t���?���%��k��[�Bt����܆��x�SN�������^.vC�IEmZ���k��D�����-�@:���
���:��<k4���� ����mW�Ωa��/�R? hQl'�?�u:p�30�'�'"�F�?�	�F o��i���K�n��r�S�c?;�M(t�b�܁�����f��}���<�����3�$Hq�&���D��0�Tkc�I�Z�Ĝn�ݯX]J��	l_������=�<�V�_���I�y>	�;l�"Qa��~^��N��e����顉��|�1��`�~p�u8��$�pg5YEcy�������LH�t�,q>�9��ޜ
�������Es���b���(p
g�uYW�\�h���b]�:���Y�p	m��5�����85C?��~�2���A��4H����S6*mGӫ�F���h�(\��� ̛q[�{��/�.WU�H���σ�5܇��x�,i�x���p�ڊ�bLK�C��de�M>B��KN�M��`��++D�<�p#:��n�RW�g�Wh��vI|q������8�Ǉ�bY����~�7�(���euk���D�B_pu�|�$!x�t��6��r�x�vxU>J���ǚ�*���:�b�A�1�B���Il�.%vm[B>xU=
{EH_����h��>�eqC2��Rn�7��7,�b�1�4��qs���g��fSbl��[>g�v6�`<kH�K�a[�)��!��}������/-�D,�a؏�b~� ���:�x~�����ނD� �g�����ʑ��-p5���C%T���&8�=���uV��gHu�W[�C,P��b�N�*k �}[�ڦ��A���o�����+�%;�_�;��<%��x����-H`�8|�`l��¢��d�v!ݥ��	�-�R�Т/�[�^I�G�u	"0̟!�9���f:�G�ڸ8�eЕ��ߐJ�ݓ��shb�8��"�mJc�)�U?��rT�_��=���<ٷ�WDE�Ȳ��2��;j�S�?D@ƚ�eǶv�+*�k2{�����G[Â�^3��]h*��S~0|�D��w��U�,����`q����e����%�s�����X�s��h�ܣ�bLCQ���*����
EJL����h]�6 0��e~H*[�Z��P��f���Н��N0�j��P""��n�7��ۨk�=y���%\�v��d�-$�{���ӯ��u܄H�/=�w��z��4^0�)��/;G	��vٙGD�0%
)fP �����Ȧ�S��/o �:L�)cq�p��V��J��a�"����,eZ���'E@���1�K�u���:�^�ձ���NDv4����MH6J�ex#�-ɷ����1��n*7g�L4�y?�Hj�b!���2��ոd�9e�j|{���ؙ��1{�yv;��n����r�UA�$\!c;}`#��gfo>�5�/�g�X������;1��#���k�Gw��%��U�WV�-stL�P�@���C��'3���c���L�	����z�I��N����*�#>�MY/��Η�4��_&K8�b��>"�6�I��\���0BU��;%�r�:�C��0�޽pF{e�?5�*�?�y]VE�����Th�A�P�������n^x ���^x����h]��4�Z������F^�K�ZK�]�Y^�#*δ[Ef�W�,N�pfݘ�7�
�I�*?��X첃�e��nI��{�c����������/W_:c-�`��WBP�5������-+!��VJ�?�5�t�y(ᄪX5,AC�����&�Lasf����<�s��<��	N�JY�\w�	QǗ
�6Q���ښ��q�4��*�b�b�g�J����x���S/W詳�M��](x����b	$3&��S	�x<]�n�д3Юpl�-�؂a���j�pgO�`Ȗ)1���!�L�䖡�E��s.��y�������;3\���,���_<<Ά�@IF�b|jR�N~��9#�B�CR������9�S5_�=�hJ+��y�N�M!&zX|�{�|VD�ck�O�	��������;-1���gb^U>9'��Eh�'b��������p��x�6�r�2@�ڥ/��\��;K�i�E����d�:��f\�[H��U׹k� �HvޯLr6uZ$o��Cؼ��ۦTd[�<A�<G�Y�BGBR�������c����|	g����N"NH�:[0s�۠8��Ֆ��y��7����z��D��X��ǯ�]�	���&�%8�?�Կvj� ���+Ϯ�pY�=�f'2����@-�i�{8��SW�]�V�J��<D���W��j��؇M�H%����_5c��|�B,��[M���>��%$L���*NҭÖ�'�?:��͜��{T�( &�^,3\[�v����|�������:ϋ�k���Kol�,��Ov�����+8w������gW��0o�!�lهW�/�)vo5�m"$���Fh�H)>(E���;�R�]��Zl�6��у�2�b���tX�mfE�?��\M�SSO24�M�=�Sƴ�?<�E2-�I�KW����B��u����k�Ga�>�M��(�N�Ƕ��;G�,m^G
ؑk��y�	��IU!tK�d�W���Y�#(n�P��'�rH0��\0{5,`����}��[q:@-��Ǭة��e� ؓM��k��%�>�kn�-�dV�C���C����yJM0��.��z�2�qŔBO���K��J%4Giҙ���J S�
�CB٪�SMp�������I��4�'�HA��!$z/=]�0(���vUb#��Mexu2��u��I8$Q�GA&���C�`D�UBr�S2�9��.������E�8tuu	�N�8��:�QǨYweg�J���M�K�@|{ڟ�?e�怓�����|!��+����,ץ�TW�ak�5���݃�!�c���������^SL�s+�ȌI�V%�I�d�]�&�3�.�qR(	���F��y}H	]w�;)h���i}MuU��.�1�R_&j%
9b�q�0
i$|j`��L�ȡ4��1����l�⌶@�i}и��S��E�7��7yh�8̳\���ED��1���qva��WV� �������������a�����p�Yъ�#��٥ȅl�@X:/vH�x�l ��@O'&c�"n�=s�2��ΰ^ZDI�ћCU����䗏��^�4u�f~��0~��X���LJ<UFR��zB��ȏ��K�/-G!ǋ�:e^k���hQb��T��gޑ^ ,�W�@�������5Y�q�`-�|-�h��qr:��(*WG�H�i[yW������=�m3vXj9��@���~eREm3�Q�����6hIJ��U�`#3ze'�'���nG�Q-A7��  $wq��{-@���u�GW�q��Y���	��ސ�/O�:O"����rin��~�u����R��%z�'�R�m���ܷݰF_��B��@aY�mH^��B�42Ҕ4�*�G�Թy'*�&�>�W�Z��6�,E��ꑿ����g�ԉ���Z41$��-72.|j2���q6�����]@y�<�s����q�-��j`*O ����	'��M
h�ɳ#Ph��s��5_���:�o�R1tyu���8�;��7IC8)%L�B�[Q��E�#�ԮV��l�5w�mv�.K�'�ݓ��|<�z3���{���z}�'�kEod ��L�F���df���~{5z�b���Y��B�RI��N&���j��)[8�?�&I������B��.Iϊ��Vh�W^�^>�-xHm�� �L��_���Ys9�P���"�Z�3�����#�T��07���}w�ѿ�����:���|�$�����I�b�-����t
�o�x�l�T�o��&3Jx�&�%���F�Ul� ��S��}�7��&+����[�8P�16��2!�x�H���|�W��rЈT��}R"��b�-�S�R��ё��2���@�U$�ZzD2ӫ���a�=@Q�G�,4s�o7�O ��_3�/*Dq���8��5ei��A+~���TQlD������i�[B�Ni�Ӫ`�M�6��0�S~�o��/_3�ZΦһ����*|��-�/�<##��_�q�Z��9g�?f�e���1�-����m|&q0��p���nl8�lGhx�r��}6T�����km�y���8 Q.yGD�����j}��{��R�j�~.����$�z:XfA:x$q<p&#�ʧ�ů�U���,�#m�K�o���ZS� ^��;�ܸ�ؖ���V��h��|�����+�u�_m�8y�f"Vx­���N/�|^?�й`�&�N��l}�ko�iٝ$�Q��������!&��r8��/i��3!�ƭ�y�+����L�9�%6��lL����T�䂞��~��m6��m��l�/������[?�b#��i�߹���Xg����s�D� �w��&�ɾ��g6#ߨ�I�a�6L�5��՚���: �E��E)�-i������� ��i0	x1��U��|b�A�?7`�2�	̆�[�X_a��.�mOM��K�s�\ۚ�^�X�<��q��m�h*�Ŏ<v*�D��Y&���Q3H�
��k�©�A��xQȟ��z��n����z��+}�$Z+_F4�R�V��^���^!4��a��)RYM,��� n�����.���С�ʶO�=��r����Z��QG����Ӿ������b1�#Vxt���4^p6|�������	���*��ב�M��h�B���q;f��``O�~*G�ՙ��Czw�pY_H���ϛoH�JF����h��(i�)��D���H҆nl��#��<:�N����}f��O;�:�5f@0�P�P7�gL�L��p����k�gb֔�"C�9��$��9�ڤ��h���]��ை,�j��%�3NKS��⚁1��ᰞZԥ��{U��*9�/m�Ƿ�g�##\�1�i��E_�o�)�q�۹�tk�UT2XMԯW��^r�yT���(J"�et���:�A��fE�_�󻒾.ſ�=��^_3Fy�%TN,�q2��b��z�$�1XV�7��8a�fx����f٣KDU'D�0��L{d�����^M�1��t�����+0cFL��6��Gj$�KK�����[��>��q��.�.�'H��i&L~40�x|�l+�v�2̸���{��&�es�ʋ%�������c����-�m�D����r��\�-��W�e&5Lc��O~v���"��q��x�3��benFl1#��m���ÂJ��@�����߹�S:P���>�A��j6�{Q�����X�#Y���iG�2�@�j�C��l[`� ��F�����ji�S�d$��"�7.fmm��t�Ox�-���^V+��Y}���8�2msWwD遲�	n��J0y�<iu���-�5���+�M-������A�%�Vo�?4S��9E��_=��2:�����t�����$3L�Pfal�����RW���S� ��`}�6@��$����VI����~̉2��B�v(b�l1�o������� �Zf-��J�Б���E�׹��z�gO��"p���_��w8�F����z�zZ|Ow"�,�!�X��G��T��4&Z�4dޣ�]����������0�Rc�yƦ��Gԛ�Њ5ć��ں��L%f|ґ�M��exh!j�x}a�Yc]3W5��a|�*��9�bh�_��f��F�ӽ�D�Z���:�E	�l;(�Z_��{�
�R~��������k8�|Я���<#C�O����s~Jr �4{o���^����b~ϱ��_'�ےң�|ì"�G�w��%s�:#����D4����2EVg���'��#��WI��|��ۜ�Ό@�*���lpo ��3"Gbn*b��a�͒e:)��J���e�'�+�Ѻ�2�9Q�|Ɖg����cf�ڒ��n�
�:��hd�٦E�<J�RCq-��A�փE
:��Ӯ��2f�@�8�aEVA96m��r���诡���M�$���-eW�_��+�I?�!!�i��O�'� ca��}�	m�.f�v�LA�T1U�%jr:M��u{�g1������v�=�g'El�	<9k@=���?�F��]�B���u�^�Z�7�wC����ɿ�-$�Y�7j9�������K�(�j5����^�ε�i�?�P}��S��Ca��X���,��(�����9�h����,F��K���2\�����r���K�n�G�8���-^Z���$*
#�����Z5I'q�ށ>��!�|8��vqZa��3�h#1�!G04OŊ��grl����˄�|v�c����PG�9zT F�Λ����-
$Du����}����p�kpo���<9�	�h!
��u�WB?&��D�$I���Þl��fߙ'Z��|�Yp��Fx)l���v��.�,\�"{yJ���f*�\�����o޵��#���]~O�h�ںCp
�n�b�G���q��B��*�iHK*�ܴ!�|-��&���^�ŒL��<�s��B]���Y�:��{��xa�}�E0�ڝ��I�V)���h�HQ8���'D�y_^q�خ�z�55�-�|�`����z���k��i�v�����C�e��e+��d���Zl)7|ˢQ����Ǝ��D��-�2β�p��<�K�/��8[�_�:�"#.'��Rڞ�:���D2�מ���J|w�J��*�������ڃ#o�T�ѻ�B�C)������`���O�N�A+�zjz*\�iI3Ij(�+��2���S��*N�����&�b�%6��$m��4��Ò�e�~������K����J�n��s����FT/�-D'�Zb��͑��K�H%^Q��g����^��l%��R�_1�U������k�,�
,gT�B�
��ڮ�bHd��B��]��,%������p����3 �ֵr:	?�2����J	N�]�C&1���&����ơ���4�o°�ng/�P^�+��B���Qa|����TN�Z���������|��A�-�D%rd��x̽w�i7�B���]45\#kyo��	9�[~J���UELj����~_�۸���΀'{W˔�)5X��1�܀q�?��k�$����(C؞;OQ�\XQ;�UR��[YCJ���������LN���3,����i
�n
I*WL��p���c��2aEsd@���׽J�ð�P�����~ ������a�(��def�Ԓ�AVS����$@_ww'�u�D�z{��`AҞA<���y���mŷ���G�=��a.�����O��:�_�9�!�2V}�+�k�c9HB�t��Ze{Gdi�z&�B��D@slwu9x��k�����uj�s��}8�9�Cg�u,�;O�yJ�����?�ζ�N�`�12b��iD�Y��y6�T�D1�>��Bg�%��v�������uVb� 
��c�㕾6��d79��q��M��8�۵�W��^$:�5�{�,�	E�</���I"Pk�Ų��4*�c?�N��b �wD"��j{,MU�r�9�z�ȫ��c���ٙ�6j�WD;wW^�����9�-T�2K�4z��Dϳ�������B�;�:�+��,�j�ڼ�Y�ox����ǔ�mu�p��`�@������u(��Ӌ]�C=�LR�Z�ް����L8����z���M1������!o�]��Y�&	�HrH�"36�n�������
ށ���9,�(��?�g"�s�v+�E��aJ$���Ö۽������}�'t�L�<T�ғ!������E�	` ��7u!z�\ɜ���`��S�Ъ�d���� �EӉ��NȘ|�_M�L�D�U���"�	�/:^Ǆ�0N�;�=�<h��� ��ZQ$�zSƙk�XOZ�G��xE8�2��ɠ▟�f�WJ����w�k�~X����3�m�$����ac�98VkS��������$��xTM6G�	$q��y�[���itČ,��wl�a8�f����H�`���Mn��Y�}���K��>����1�@�>�ң��������ąY	��k�Iפu���o!�̎�e]Y��H��D �������������4�s<)��樲���7' `��=����U�dO�͏H�o�����I�#P��-{#^}�M�v�t̡���ܱ(����d��R����y.�F9l�}�?%�/HG/�̯8�G�w�M�O���:�)=��X2�-�����A[HI�w���~�����F��ʎE�K\ߐ@�-�������8��	��z;�=K}��7T�:��j�yz��nb�n�H�{F���2h}J)E���/����4���{ܯ 鬒�Pj��z���ۥe���U�/�,R�,kH��X:{R�:l�JAۚ��8&��{�y�]�p5|�K��Pw��[�{u�1A��J
^�M3P�@)C�EI«W�q�����85�54�Rq 	y��n�J��*���-:�:S~�l6�������OQ�ْ�,lb��@�{��F-�\�	nͩo$�'D,xdKR.�J�
Ri��`tOh�&	�)@<
�X�uFeQ�sʆ#��(�/Ⱦ���\`$z�yI�U�l�^���A9�a|8���l:%��@&�/v�"C[p��,�[�����?-.�ӫe�:��n#�rO��0:��rH&,m��Q�����д>,�#S�6{�~Y<K���UX&��C~W=C����c����� �IBc�<u,kg��᫁�*�xX'+A_,M���A��ș��9IW�ȼ( ��m�.���(u!.�u��������i�>W*D���B¬u�0� g�ߠ��t
Eߨ��ҫ&L�=�������ë�q$���gN����2u�cCC P�l������♡��P���a��Һ�����j��)}v�ɍ�l�g��5K���T�I=GC��yL�|@�0g<?;+?�?�p�~�O��������هX�gT�)��	+��G�YP�ւ�aVX���2��`���'�}�=(��_�T]�a3M��w6/tkw#��`=v�7��ͨ�K����m�t'�ו8�>��ꮎ/����f��D2C�ΌM1���\�׆�S8D��P7!���'<����$ܸ�ק4�-7nu����S(�`��.Fd�����k�s��)�[��|ಈ�@��3���Iۖ�3,wP)�er��l��Sh���V��N�eKU$EӋ�;��ŀU��<���U�1x�w�Fgz��%�vmSQ���iY~��uIٌ�`���L�ٌ� SQB��2�����F�T���p�������2�~�W&eI�+^��inh)�:�E�AV�}h�63r�p�zf�q:�q�#'��6RCH�(0��#��Á	�d�oz��-�E�w�ȸ\�ȡZ5�c��w�dU��|�I�5v��\�v�� � �-D�E,=cC�i���6��'2Qq>L j&$K�:w3lٹ^��gO�u��KD��'��(5QKWē�*�?��}Si��@ϟ�Ŏ��O�d��2�b�$�w{O��8Z'ǥ<x1#��&Or��\�xă,��6F��38�^��J���C��ݒ5k��(^����Pi��� ˒.�h	9�~��k���M�5G�1�0���C>j�*A�a�WZީ�'�О����u�R;Se��5�~^;2��%�-{��e�.]�|8��`8��xr3�[?M� ^֘��uy�k�#-�T�a|ɗH�Y;$�3�(uvҏ�\���-K�~��͟�0\ ;9� ��*3��;��k�����pi�7�˟����N�F9��U����5���|�7��$s}_\s)�&�l�sm^;#{X༐�U�St��i��NMA}r�|��^s�r-햬���I��a�x^�GY��ђP{���=�����Y���^+�]Ϩ9YO�n8�رA6���1�l�p]�����D*J���9|4��D�h���9c��rW9��Y�ִ�L�������*.f�Y�-�X��X��_��{��ug�N�h�X�ȃ�׏�+�����R�s����2UQ��y2b��Xm�D��+�,sJ����!
�m��I�n8��s%,%E@�c����"�e�D`X@��
P<�X�����~�j(9�������n@� �ε�`�&U��*uߜ��G��=ү�#у����6+�f�}��?�{|���is�!2)IU��&�es�H�&6�˱o����fL6m���T�?#��dS���=V�@N�&>@8�`%��~2-w��w��#��|,Q��0�{�x�O��\#f���A��C��˭XdP�Vd.�V���=�
^��%�QQ�%��$�2������w�+�r��.ِ��e�j?�Rh8���`�{]��1�D�bbڜ�z���/2!�N�J�g�7��/��D�B�Ee�Gm�W�j��N�VNI��Z�!��� f
#v��\��Q����o6N@�Z�U��3wT�"� ��ND\>Q���k 6)-�/��j��Za'��tQA�H�_5��h'}�K d�亠��x
H�� ��]C��3�٪�XC�����'�c����|=�^�m���7�S�&�^o��(�d��_n�P���>>�,ș�4P>M��V���E��ν��k���M^�����T<�e�A�2w}�3��i��C�-,e����ԟ$��Z �cA~V0R]�^��LS��r
����V
�l��{tV��hS^`��u��'�	��0�<��<s`S�2w��륎7�"���8�i�Q�)$��m�f��E{�hc�]3�G3}��8
iy�����Ӻ�N�����|��)�.������S29���w���䑥��p� 9}b$���Ț�$�{�.|��=����]�����]�h�1K��cnџ۞��z�J�3�0tr��F�*h$� s��;=-�YRY䔧�8�����:D� a��SG<k�MfT��|�%�^C��!H�öv9M��s]��^G�� �ڛ��X�(��V��V�C�ǟɻ�����w��ZMe]��Xd ��h�a�!!�<6��S��6�;Nt��2J ���t�����D�)t���#K�8Ys&V-e��.��X=�E��u��\,O:�\!��t�s��CjW��u�h8J�D�-�K�dt'�"�QaR�w�Ϟ�aމ�:��]�M�N_��/��*#f%��g�A����O}��'�E�T3����a}8jQ��:vsS���E8�������L&��C�k-'��,J�p��1`�?��dk�m������%kh�Fq�6� �Wr1�+(A�!5�:��g?����ϖ��n%�/`�w�L���a�J���l�� `�&��)�:��&{f?Oj!�;:{�%4_=0�s��o�4) �+Ǣ4I�����W�CI.�L�M�*
���d�Y����j�w�ë@����A]ڍr���I���.��
�q\2�5ʤ.{�Wg��D������c����{����%�QM�'/8�^�~��T/�")�����>�zg[�OݣФ{�b�m��I�v�I�Y�.G�3=`.sث���V�l���IV�����~�!0��gQ��O�p�*���Y}��&�'��.q��&��y#�<|�y��.��i��(��{<8��w��<WF�-{�NP�����P�(�R%��ub��;�C�2�К�����cg����'X��7w�(��`4�l,�e� Bֺ��#��j�L������ӕ����qY����e����b��6�n ���#�kn���2lZK���,j2zQ"�u�ˮ+rT�)31M�_,ruSN0W���E�U���L�[EȷFɰɁ�y!�(��&��DD��Q�*l�k�WU�匢� 6�x�o��4��9����Dc.�&'���T�U���g��i�u����~�$�ȏy5���G�2Ϋ%�3C�m�!<߭/��z���f
��4��|�@�L=�M꬏&�v�X�%�c�^��$/�7{}��9YO�:aF������{�@x�s-��A��q����b��9��~��;�%�����N��Y�P�P�ڴ��e0x+�n�eЉ�h��;ǌe��ٺ�K�VO�ĺ�Љ�ޢ^Ōy�<�Z�������Q��˻�^$���N�6�J��s]
�$�e�^�Ђ����!\0�a ���m���[�����8�q�Rn��|��s�/0��͕`KS߃�$f.�8˹ۜpM)����P;7HUfHXcL�J3�8��1� fB�r�R:	�d޲��	'f�r�o,j/����R������gkC�f�V	A"�g�kC6_���Y�����	zr��s��e��떞VA�޲:���r�}j�/��w� A��a�L�MU*� +}�Q����ܯߺp
�S�}ep�5?b\�V���O��~�p�0$4��0]��zz�yo7s�b:Z�dRAV4�ìl�Yx����x�0f�5���'Ʊ���h�J�������<�'�u*��[g@
��O??�&A��k$h�[�~��j�9�W�p��'h���O�i(#^��-"�!�''~�TΝ�� �÷�����*�]I��TC�����s�������5��R*�ލ9�����Sߪ�n�
0Q^,���5����5My��tF5`ЍAnB�ex�%��Z�����#�$���E���b{�G��Wpf�n]��`��/G���ށ��Zaﺟk�g�g�e�����d�[f��fM�e�'Y���������5�s��)T�� p���V�v,��
@�I,�n�hv��e�q��������=>Ӓ ��K��Dt�镣�y,T9<4.̯X�Hb�)��E|��ǄlRee`=�	xӁ��]< ��l싯){d�rT�by��?$��W�΀��1�䝻]��n����3�����=�������� �S�����?�B��Wg��@f}���{�{"�}��rV	����w���PŹ/ok� X �f���s��B���#��	�R�8=�_b �uSRn�I��L�j��t���]Ճ+��3�G����v�ung`�Z� �
�C�gO��­�`�
�/��I�+��,�P���l��,S�~��	�Ɏj"w�0i_W�Ej��� �b�3߈�gq��l����Zb`� 5����4i�8�S�r?���X�ڀ���k��͍���=,�/j}3��J#hi}|����ޟ>��p��/^�&cdA`y���1�y�I^&�v��U�]<y��4�F��5�ͷ� ������N��A�"��]�R �;� yX?��'����*�9O�4��&?bi4m�&�YK3B��N21�/�a�3��Yd�2��:k�}>npc2]��H��4���`��!�.Z����V�oޅvM�����V�{B�����k���gتGt?��Ш�� '���Jߡ!�eEu*��;Xz�j[�V��r�X�Q�KE������ E��I��?�����K�� E.E�I�����V,斘�PX�A�|E�l�y�=:=`�"��~��l;�ɀ !�=�m?���w)�9m���=GPG�7��"�g�=�£���ٙYS���8%��(Q��l��� ��w�N�[��T ��x��O(��˭%��M̤�a0�a�|��G�������2��*F���mVp�\���;T"i>��D Wʘ�4O�h<E;��r0۾�O�a�����_q�(��a@|c`8�^����Bk��m�+;�^�f�5��5��#��}�����Kl���Nם�"4�X �p�]R�u�D`�����װ�2g$^�}x�!����{x��"<��ƃ���&$W�1���֑��P?*��o�8+ Ao�xÇR�ΜP�O�&ϱ����E���uW�"m�}�/��D̗h�Tyl���^5!���;A{�y���We#W��X�av�l�ˮ�Z<5�V΂��>k�װ����A�5@d;hS��o �~�!d*�R�F*ͭR$s_d>weCR<��!�g�2�K�}���ż����BX��uQ��q\Ur���'_.���MR!�,fa�C���5��Tm�JO<M�[z~�*�Ѩ3�8O;�$U�B�4&�)�#�t�NC*��Q^�b��Oeꁵݓ�#�G�5?�:V�m�/��3v�t;�txp\��9+}��CP�NOc�~);`=G¹kzh�RsM��LTe}��v�g7�C�2�ʲ���D���,"��Jԏ�T�̄O�w�ܱ5�8Ỿb����Ѥ�2����Κ$�!�7����
\Ջ�9��'ʍt��$���;3Ped��M>�3�(L�d(_����e���4CMɋ�{^�>GwN���:Gp�J�F���Ж����T��:Z�7#�Y��kS����m��f�M���%uD��	�O~|@��U[�?�>�4���"�Qq���s=P�ɦ�#3R^��&�#��-��I2���i�3�ܶ(?�tG�&g�̐�G�RΡH�2�5:B�H\�-=?���Q�+��R�ŎԵ��ä��?Ev'�*w����I���c� 7�L_y�M�%<^�R<�o�O����r��� �}q�#/C��o�ft�I}�3�ᝫU��t1P�gc8m��Y�M#!�pPMx�0�Y�x!p,O��E�|Y���5`���"��8 !M,��J��5�����ހ��e3�Ǚݒ��#�O�GI��[<��A_ĩ�s)���C]�Ǣg�Ƴc��VD|�MQ�%!ss��]g�����I�g��4�����N����8�>��oV�/a��I �e=��q�v4uB�WEƾ��~�9%Eh�L�*H��B���K�n�n�ߝ�={Po;i܂���n��0�\�&aDD�vb�Q�JhG�'∰$}��v[^��i���X��d~��5�\ѯ�C�e�&��?d�V��#�ΡD9d���ː�鄍O���T{O&SdI�_�,�Tm��R =_�*xl��h�%A���T�ϐ��yd�W�;��e!�p��)'���w�1^j�Zoi�gR��޴?�Ӗ2&(��w�J�ɿ��Y!q�)���Bmߘ1�h�B��|z���+Ny��`H�`�JѪ�x��̌>�&3��.w�~�vWR"�[������"���[�����)��vW�d�9�A+�"ۺo�P�1�ZU~��O�t�n���4��;z�Ωq�K�~H@>8x�|�ѕ%�K��8��<
GM��%ebYfB�}:3<,��ۓ.�箨Z|���45���KfYS�+c���~I҃~���f_�A���G��2j>On�����D3F@��}�ؔ_%5�*:PzN��=A0Y����y6/:RO�^�f!U�o��;v��U��c?���V�z�C�P���K�Z�����&�� >��g���[E=2Z�L�ގ�"������PX����>��U���K�[~��S�t��rk�D$X��Ըf:T���� �1L��+ݛ�#7�e'��V���7m��!�X��98���ނ� �׍�`nE�?�=�37-�7n���	�TS�y����*�'�"�bH?8BH+�ذv-�>� &w�ި��}�ǧ�989p��S�ΰcbF�{�JT���f\�5���2��M��j����3��	j�T�K=�x��**3���T2\��i$W�6��ҽ��K�cJ�C-հ\���bxo���|
��μګ~ٸ�t�����x�ĭ���յG�t@���`a"!�6BL�s[���|�
�Ϲwŷ������qd�����Z��\��ȚL#�'�j갿o�T�s���F�U��(ô� ���#�pt��@������js�qg_lKT�[G��S�E�@\�YD09C����#�`����4��fY�2��������e5�d��X��j��np���I��	K�ڿ�>�C�����"����a�M�PE�[f�t6ۢ�c���;y�Zr�!��aL��������f�;�``�.cu'����_�['�2�c}-��;�o���%a��jw�/�=&��HeIũ|
V�!��f����2<���m�}cO�5���ަ=p�8��+G{��d��/,��}�J����{��p�L�|�8A����y".���rV�QA�a����D�|�G61�
�LR���A�(.�"��S�"\�M!l�V�ڶ*ʨ�.�1L�v_�'�OIC)��$FvpY����_��V�l�wR?��q���= �~!���fl�m�=P��4���`v0��p@ėk�B�!3�o>6imm�״�X�m� :�g��|Ց���t��DՃ@Yc�ָ��x6������������`�߮:�sjrn8��w�g��=��{��el&5���I�3��;{@c��Ф`��(c<4�KHygY� 3��~|$st
�B��r�D~>f��!ib,���qK�G�H	g*�7@���Hÿݘ}⿺a���y`�D�i�i �liN��M��s�S�b����Jɦm�k��:>_��U��_/��1%p�K �:V�Fq� ZG����X6	�u�2g��0�׹eN��y���N&,&�ܦ ��\9�����2��l>�3C�������K�Δ�c��v����(>߉&�W[<���1��?��^K�����t�����������O�R�.1�d��ؐ ��O�\#�q���+��Wu	�Ɖ}uuN���r��c-{�*�qڜ%���ޣ����Ժ�(#H�W�>˛��_k[/����z�j��>>�G��#P1X`�N�e@��F���)\�;Bb�nﲉ���k3��LP"�����V2n�5ʹs8��⋑����G٤ނ7�c�4�''�Û����g#5������Ǖ�yqPe�vqkm���K.�L&K�C���_��*�5̮��ύO�B�X96��
Ԩ� N`��U$E�����.��8bz@����ɂi��X�x�� Pޡ�2F�uV����#e���u%����Q�Xm�K[��0&{�����<�'�g�od���u4oB������\Ð�W�Jh�K/Q�b�غg�'.&C"����$gc�$F
I��U�,��n���r&�g�mV0A�Y�w�̾p��[B�H����۸e�q ���柙N��ꅷ�ȏr}�G޿9OCZ`z�2r�B���N���\��E��y2��z�5B��DW�Tt�9qzX ��6��~_�b�������Va"������N�|���׀T�2�1o8դ"�	�GL��#��^�F`�"MԠ�W�!��05&`[Oѧˎ��*s��N�m�H�pa{��;b	�v"��ze�=�pn�j�v�U0/���P��G�e��l��p�&��jK���h�<d��5�:��N�7f#�/4�?����4ZeL\4.]An{��SW_
��/���Dx8 ��p���,޶;n�}��lI���#�����9��Y�����̘Iʩ���pSD��,������b��ne��������:��%�ᐬ���^�4BW�g�Y
�M����X�x��02@�9V�q���i���'�@d���M�;3K�,��up��u*kɺ���ej.�t�oP�9��J�R�����Ut)����s�/X҄x�AC�w9�4�rc�������_2���tφ��;�K/_���Zj~0���,��5����)���Z�HBr��hW��ܨ=��-�%� �{�S7�A�W�'���u�8�p�0��Y�a7zS���������[I�4u�&p�ԖC�QJ���%�l �/sY-~�q�U����$\B��n��������6�:>�a0�C\|uY����?ǻu�&i��6��n�|QY��x���޻����yc#�HәC=��m.{�^h)l�K����v0�&����yv�Շ�)�,�QL�J��MC�"偏��zw\����#�ऻ�%�V۲
jo';.�T�d 	���7���X���+�Q_>B�aJ-9@�r_� 5q��E��~ߖ����uW�D|?϶�6�b��6���=Ke���E�<��7�ʕ�R�������@Il=�|)#�.{���6��Mi���G�R�n���&��p�����čp�$t4��N-��A��y���S���������K��";�M�9��������o�C��� �����)�@0EX�܀1M~���ꇗ~�ǅr����+�UI��O��#2�Ϝ�)�#����LcR�:��7JH�uҍe7 .����S�&/�P�꾰^i��F�������\0�u�V<�\���w��̜�4�j�� 
���+3�nP�)�ݫO��ʃϘ6�>p�㰧u��vI�K�G��+����{,֚)�t���fE����=A(��2���[�̭����3�=�m����t�����k�(�.k1��[x��p�4�m�{���xMƑ.IGFSƂ ���铧N_f�t�%�1�����s���Al���lE��r-F��c��C�jiX�J�
����>�˶I�	Ff��Ω�@Q]�y~'�����?_���x��X�3��Q_mU�3;Ht������m�@����v�4��NO�{�~G�`k���,��v5��Q
�5z ��љ���6�؀���i2mo}~��z�!�>t0e)���7�(�����E��ԇ)c�5B+hCf��/�~k=�T�t{"��BǃGc�a@w1X���B&b����}����P��4$�<��L[~Bz���+���L\mҙmi�ӨУ&�_2���=�-8������t�F`��;�#��{�@s�d91�
H���hX�j@��p�'�)�I~�՟�[=��}���p��H�"+�gl�%�l[&�8$�A�u_�ڠ����*�V���!~�񶾞��c2��+��	}vp`�_H\���_
VW|T����6�j�[�f �k���Ut���'~��^mcͿT�A��Ɂ��@��0'��	;�֍�<��JP��G<���g-�s�]��7��XR?*k�Wė�M3�[-Ƿ|?����Rb�v��o���3H�k�p���4&h��R���b�gT��^gSR�����V6����7E�!��wc̐�h��A����R�� Ң�7SJ���e�Ո>��A{��b��k��h1cl�hF��:� -�F��{fɝ[L�v���Q�/�b�j��m�����;K������bSc3H��lf���3�$���ɷ��O]�!L�(8����Vs̠��AK���)�o��h��ꪉe=������qˆr\���+]�-L���`��ԃ�O� n40���h��Y�6�O��W.`9^���.�+�䄿蘬 �M-��*������9�ag	V�Z�8��w��S����]ԁ���EN�����1��m.��j��f����Gd̃����H�JOz~��[ʩ�J� c�#
� z;�[>�r�d���qױ〮�ت�wA��z l&���04vBd*R�������6�|Y��8�S*�q� i�ɚ��97J�8�W�WD�>}@��j�8K�(�����x4|�/���NE�6���ݢ@����
Q7h=���.��yTv([·���t���?6DY6'

�jIG#Ԓ��g@ sYy	}��"p/���y��1��n3��@p�EQL��l��MSg�:��\R��&T4�U2k��Ҿ=�V�f�gk�A�[ �;*/�-p�U�?�Aw�
��s�YU�������v\A�I�d�4}\�1���u�7���?S	��^I3hۨ/2�1�C$%ۥܟ���j���䕁��=�S3o�BMi���T&P4��5��x^5��u��i԰c��<!u�=��"e�:���1�b5�ݝ��
ۭ�X{A�[Lɗ�U�p�:Y9hF3=�Z2n��FZ�e�o�xF��Һ�����x���NȬ��_1���l�p9���(��|�x�����K\X�,S�3��3�b��(��2A���L+��i%M	�/�ܬ<�oJ~����K-bO݅�r��{�8V��>y��K��ʐ�[C�p���\Ts�� ��H�`��Ґ5���r=s���Pa���J�
�9�脘~	۟�=�-|>�h7��Ҳ�[�HOˮ���9�
��6ю�Ӱ;[d�Q�!�UDV��j7��V��R:P�8i(m:���C���旽�Q%��ۢ٪��h�V�g�N�$LH���`6Q��h�_�uS`*��ȑ�+aZ
,�)��j��v��3�	�����p���X]R��Cxb[9�rg�Ca-C�K��H�屩�P�y��30��0f^H.���x#;u��vzf�j��,�&�����3Q�B$].Yzpρs���"�M��4�x�\=`��a���]��5����]/e���D��)*�d�~nZPݖ�By�΍��K|���kg���Q;���}Am��j���ӎ��Wfc!�D�ڞ�Cd	�K�kT�>]�GwRR�(����^fW�<~���hl�V�d���5��*�E/j���d�����p����1ŦW+�"�r�#.Mb��Tp�쬀kc�S�Uzbp�F=�G0w�ls:#�8��K���a3}��+��U�a�n�L&�VAgB��_*k2l�S$��>�k�h"�<
%�W9�z�C;u��g��?"�>ܖ,���R5��h�H��: �p�Z�AjLN�����Յ�^=��H%�Q��f�U���_f����7�n+���}���3�����9�4A�yC[?Y��W H*�Y>,>yJ���Hxw�s�{l+ �s%x*Ջ�c�]�q������ZeH����pe����B��%4�*H�7�����J�� �Ԋ ]D�g{P����gJj	�|%�6Q`�!�]b�|�ΐF>ca �!����z��Q2��e,0o��/���A|}z%}�@�[xy}Q_2��J��§��P����Q���\qop�7E�+�j��_���FMA�H�D���xrԐ��4'Q���d�ZtEω��ݙc�h+��0+�T�Sz7��W�:��V3	��R�������_K�9��L����4�^����mӔ�hk���Jvզޠ�Qn�5�&�[WZ _��8�y`	�.��gh󏇫JS�� ���Cx	��G��� /��_�$�7����1?y 7D �Dsy�W�A7k(%��qu�J���i9��y5�w�@(/�{Q�Bg@p��/��|����?��E�]�l^�ڇW�/���FV��(rhi|r�7�s��t�Z�f ��",����J�FN�`R��^ܿ���y`��c�`U�I&��������������0yi+��{4��jIY���^�E� a���ʘL	�fP�f�p@�ΐ�E���E��Ojk,�J�!q}#����?�e�h@��*MM{K�^��|N��X���
�V�[T��t}Qb�m>�qƁ[����eM����M	"�JHS�K7��5X>��2�x�{ �~�c���Ro��]M�P��L-:�qF�v_��"5[�>������~���v�'l�zb��R��E+·�K��<�`gZG�3cI]T��uG��&�zY%=Ҡ��r�#<�:����d�5"�U��>0��r-;��6+.�������@ge�c#�fЂT'g��9h[!m
в�&@��ڰ�|���s;ֽ��~�����e�Y��,I�����:�kg4��s*��nO�x���)ݟ"[r$��5NXjٯ�n��k��" ��dX��]��_�0�l�`[�*��.|���E��\�{̈,�M6���eZXm��y���?�;8��A�san�*zO�I�ۊ6bP��qʜ����Ë�A!� �0y�&��ٸւF�ʐ���f�4����8�,�_ui�#R��I�p2��~ATN�\S�p��X�<�	���;W��vz��ݕ+����{���1�v�1���;	Ϙ���s��<����47�ÀT��φ]4|�!F_S��I�c���K�(,��$�R�Y�����#�0��})�VU;���a4o�7Y$:1,�.kwZeދ��`Jxm�)�����(��"���y��Bi�d�~Q.Y���6汨�*�gF�`+Y������'W���h��v��:���i~�B�4@B\��$�G�.�ǙH �]���~�OQ���=e:;���G��c�9ϸ��me99�PS�&�}�%>�
R��\�E���|6��)fT~e�s&:��m ok.�y�t/ف����3W���%!��v��RU$r��L�1Ik�RqR7<R_)�1��� �q�́3�Ğ����t�j�)Gٶ�2K�wQM�l�B���~[@�'
)���ù6��O4{��l��Cl��l�~�h�Ɋ$K��|�~����Q�H����v�)y�J�g�UӧH�z���48䧺�)/�"�^j��*��悜	H$�&a��ٯ����[r�1<�W��:�3�'QȆ�a��Vȷ�ShJ�6{��vH�Z����!<�x�VR���"]��%�{
�_�7P�sc��%���}γ�,��ד�9�em<��l�E+�.آ�/�)��(����>��J-K�*���\��|�N/y�*�}��� ��Q �?��zY4v��'d�}h-\
��A��$�>m����WAș��vY$T��3V��$}LůJ�dRЫs�����U.�p�u�|�'�|�|Ĳn���i~_&��^�,Eq~�,�{�%�ux;O�q��B3�Of�1ƺ���m�� g��n������	6	�~~��y� 
���ַ���gb)���O�+���l�l_r,Bb�w�t=�E��*$=]Wm+5���}e�`&7c.g�w�w�&C:�hu�e]ۂj��^��pǲt.���e��������{��
����#ڞ�^�q�T�����č�H����f�-G��rg��f�S��E�n�#�;�I����3N��p4�K;�J�d�$6�*K�s0hݓjjΟ~�����,�{�L����)F�]*�d��Ը6���1~�)�]5^x�`�~i��ݸ�0V��8YO�D9ij����NGt���QX�0|��8�hW*��Cͨ������r���\��W-,�����OVd���3&C�Lt��O%��N�I9����o^i���r�pז�,ܚ4A��4!�l�$�4ER�JCk5xԷ?�W���n�����N(�<��6��γI�x���M��ך�Q>M��z��\Z>��W["��G�c�KR��eK�A��fy�me�C�����g1Y����C�s�7U_`c	ʒ)��p��02[���F��yQ��2#�!m��L�g�3��j8#���u	j\���bB��Z�34���6�^L�ڒ-��jwn�����D-����qɞ
X���J�����J���NEOl4�����mKS~�5����I
I{w��c�3�[���vD#_})��Ɣ���t�к�?���a�ML�s���>-Z�G�;����ҕԒF�r�C�xY=!.�2�m�͈�����W�(��/�էǠ�1�
�J���J��	�o(c���hW���}Rb��kDm_	r���4	��d��=�պOF��v]�oS���烂52�b7�(��:����ǲ���H�lC��q���7�t�ד�Ϧ_��)��]{�if=�3!�}��.�=u 0y�R��G�a)P��g�M�-��/�!��)=+����sN��`�I��#��A��c~0��=�_�a3�h�G�N,q���@��T�贎h���w�L�f��ev����Lb��U[&Z���O��[N�<�^��8��6%ޣ�sʵ�#3iG�5�)��DQ̱#�Q�S��(�ٔ�D60���Z6sR��� ,�ɠPU��~]:�:S�^r��c�v�8i���W�H��� Uk&߬5-G��P҂`@#뮦��W\�h���.4�u�^w���s��_/��dv�+U���][����O�T���e��ΰ}�����rx1ժxr/�u\g�Æ��0�i�E�y��`~�b	���W���)�v>It���g^H�I^��z?E�׫<��ˬdJ�B�ń#iZ�7yC�?�#���TZ�B~�O�z��ܽe�:%OS����7A��ǘ5V+�J�(�l�~� $8p����3!��s݅$�mֈsޕr�m�^z�7x)��~s~�,v����Nw�ڹ�8�t����/I��3�;���-AVb�Sqh^G��&$�ˊb�5��'+�_F��7���Fg�"��D�3u5^,�ʗDM�|z���]
��Hφ�@�D���lf��ɥ����KvԵ�֑����^�ϱ)��FLPQ#1so�%9z��s����{�Du7ꃉ�en"B��T���-�����֧	�����͡��� П�~��K���ѹx��>j�x�m�P�k�X;%<G����QR��k�U���r�a�j���ԣr�ʉ�(�PAx�Mc�����[����>�~��Q���هc�dQ'@���I��N�ҿ��
��T���D?C��m��ˊ �wI�X����k�V�fN�1����H-y�o�~M��iA[��}~ބ�������pi"��	cw@J}�(���57q(�o�f�m_��]Z��BƇ�:ݻ��육�����_ߢ���1pO�=���2�ʆÂ.9��P$�xhS��������Szޫ�Dj�=C�4G�K)G!7�Il,�Y�rv�j�M�& ),rO!�����N�A�m!�L��5��B]��Nր�W5�5ۓ#��o<D"9��cq�B7�!�����o�l�vr�ҡ<cP�������I!�(V��>d���:�r�Zg9޸$*W��VP��(��4X����9
��]�HS�/
c>A3FYǹ�@w~L��i�6ױ��V� }\gc`�u�\���"�K���Q"_6��2r�.�޶Lʨ�Իӣ��0��_8�����̕|S�|�ܥ������U꨷�����k�%��v4�Л� #ĉ��_G��,����m���y��e�����F��p"��]
��N0�Ѧ�����$`KF D�1n=8�y�j�"Ȩ���ua����b����ښM"��Q�� �x�2�x�%�;�&Z�cvcx�M��PN(�lY�~T&~^�|�-a�2`ׂ�j��Z3��^R|"��{OI	KV�(_Vc���i���?�N? d|�w�E�c��R�E� �Q[U%@�^�s�&����բ�(@T7�
��%�>�ч���uH�!45��g����ǒ	R"�/8�G?�`L���~ �+J�/��%�DqGU� %���W S�P�4�_&��po�Ǜ[w�9������W�U��f�l��?Wd�d���C�T&�T9Cz��cӸǥ���Jl�mP��m ��٣E?��WvFz�=��u�z`"1g|��������>�&g+Tհ��P���VS�C��)K�x�����M�`[9(����.��^���������D�}N.F�s%}~�`�^�̡fh���\�lWW�ׄ�\K��,iiB��6 fT�G�2��_�)N�&�PW�&r�S�}���4�\��@t}���UV��3���m�6��l]2*|�"K_wr�6�/&:̦�)�S�R���/(I�!��at&%H\��Ԩ���ob#�|c�(���d��ڮƂ��21����}��R����{�����7m�,��qB��ۮ'*x��<[`��#�/Ր����NW��A��1A� ;��\
Ӱ�W'w{�����t��AF ��mW��0����9w3�_��~�!}����17�	C�^&�VS`�yrK�-����=_sA�PLh���S��ˇ�����ؠI�c��4���P~R5������Y�s�� �׼��W5�_�L]�<Y8�TE���������Ps��Ak�M�����cf$j�.WS�T��}Q{>O��{Ot!> xVA�����5u�}iQy�M��0��5��=�0EE6E�]�o�˒}9呑����[h��UG��~ꔤ���(e�ǻB�.��^�ܖ�.*��L�q��gmu�Rڕ����D%^qE���J��G��@A=�o���o
"�n�e#?_�r���<u�x)�-���j�{G�
Z<�0�۹�b`붆�bзqOkh���1�W�u�:¸������&켼��T�2��OqO�3��qr�!�{��ӡW6vC��!p��%��;�L>��4�6Ǟ�:�ϟ3_����Ϙ��w��و��bl�!�>aRƈ����B��U��!\@�	%�1��]L,��26nh�ә�Hx��1jB���h���^���Rk��
���[����u%���f$n_$p�CJ�K6:]1>�R�Oe腃�;�ߓB���\k�zH	�jY�����|w��F��S��I��T� ]	�o�B`�]����[_�?���Xg>�k)�=�gw��(�D�Q� �GaU�DA������J��	ZѮ�+��D��h��ސ�4���U>�P�) ǯ>���<D[p�L���b�����Q���Y��C�wy⬐O`��V�y�`sm�<����i�u�,�mH��&�7u4Ob;�5��ܢ�Wl�<�R� �.�82u��0hg��I�6�@A{(Q�Ez({�&����ڣ)��}�X�2���~eI�,7ɘ#V0�w�,����W����}�k_en(HHxr���C�nЇ�L�v�f?�g0=z���P�C�x� �N��~�Vݢ�i�5�պ���?�����+�˥	|_NUq���K�]0�Y�x�c�/
�a�U鳿"/�=���I���+���=6(�����\������j16���sz+ʢОG.��bxG��NC�?H�-��,�O�~35N}>�Q:Z�(��?ӯن�[HP�����oc8|��%^��ޛ�-���J;�yk��@�3){)�e����/[,L��Ua��޽A #��h�>н�R��Q����-�Iz�pT��l�M���Ech� ���(֤�f+BXƹ#�H9��Ʊ㿾'�D�%z�å&����W -.�Iht8��ܻи��:.�B�{���
I�'��1����@��y�Kh���%:�&� k���)'Fȋ��@��jE���[��4�8^̂�"��q��sT<Y��g_v=H^�N����7�-f�̄	�^b+q
H����1e>Dn��C�e�ۅ�g�-d�59q`�\x�d�9���>j�.������Vk�ѵ_W��@0h[�߽֤������C5��O>A�Xq`w$V�����զ7L��5�yAi���L�5�ph����맱6TB�u�^>��&�	���$2-���k���R�=WT��2��ω�gq���l��6�Wn�C�=Hc�F�l�w����qL�}��Q��i)Ң�_�	;��C�Yq/���ˑn?����V�{��~�+���p�\wc?�ʲ�D��m���Tp*���&,H� [�'qJ*Q�a�zF��I�'�g��	�D{�����l������һ�^v���)�`�``�2wir��D��z>�C��	��j��*��P$g8�9���P���p��5�V�Y�M�q�̨���<�ܡ��u��|J���' 6��Җ��C��$R{���+�\4�]lp	�l����?���NϺ�-+B�g����� q�����_$��+�7��Q�D�K�<[�2=ts��E܎'>������z�в:�If]F�=�hڃ���H����j���ƚ
�<��t��1���[��^o��S������\��ᇎT+Z�'-��z�us�F6��{�p1�%7�ƍnrx�(^/�$A<S'b����\C,�ɥ=�Ŋ W����.�{�Zc诖li";[���?���ڊ6q)�'�lAm�K|�|~e����w�����O��Q
v&U�
�?��Mщ��܂�f�$G��,qe��C��I�c:29�ň��́�3A���m�c?f�v(4*�sؾ&tl�wʴ%��f˒���"6xֿ�?n��L��Ƌ���,K#+�SCv���b|i��84���E+�a���4���VT�'Y��*�+��?v��p���t�r����}��:�L{(�D��)UR��c�C#��I������x���v-{��E��I�~S���)�\W������Ʉ��7���L���ן��.�O�\���|+�⒀J�?������P.kW=`��dJ�#�sK]�vnh�5@+/p<���\�z!����;��6��R,��b*���k�&�C]�P �ۭ#���x�E@ğJ�|8��D���w:�źSb��g˭к����J�R�YS�yz'n�I��>i��^����DA��K��� R�z!l��Z����e���*|ߊ� �>�ҩ��ڮx��w¸�����qE�<�,T��-�\�R��$������~�=:�PKT����8�w7��p�9�e����Ų�ǩ|�L�c��֪��$H�)�c2����g鮼�l.�d����w��PYI��"����t��DՆO��C�A���L`��q������l�
5-]���f��@��J�&��09��!:��"鐊s_�WiX���LaX��x��W���F�LiD�
66�?�#u[mҥՃ'иtq�Eуnf���`y�#ȭ��>�>�lXA:���W��^3J���B�K,4$���<a�r�Ev(Q��	&�3%�$�V)$�_%�1}z��]Ȥ"xM�˵rd���]9(=�K��U9�l�MWA����z��f��2wĨ�ӉZ���=kU�=˦������r�/���ֶPy&���D�3Ԑ2U
�������4������K֍�]�R/�6�VA.?�ʜ�4x;:v͙��l�;1�(�~ؔcn���ƪ!��.�5��iq�Mݦ$��˛o���Hy�GH���Wk۴���J(���'��:����+�Ђ�U3�H���铮HL61����4��O �̌����uo�.��G�m�Faf0/�M{E�P�|+Gn�{XTʹ$-g�v~��5������~,|1��o֯�I�Nˣ���Ǔ��3�����(��(�Q6�r�[�y�����A�P8BV�ᡥ�&Fr��@���o-w=x�{!�vC>��.���	n���N�	���.�h�}�"7�m��>:��Cat�A�����U'؉wL�c���#���Ir��qa}K.To3EL��Z���!�'��t�J��ۇ�|�N��������r����(���Hn�4�`V�S�O���(�M�D�V
�O,iyg����F���bA�	�B��c�]�S(�5�.�O�����'��3����UK
�;ա��,D�~����`I�g��%�`zk��A<�ښL��2���ː������e��&4�#!`c?����aEY����~ź����~�.�|0SΞ��g�������B�R��F�C��5 ՛�������i���Y��� ��B.PzO�EPU�� �D�p����D����<&�Aa�r��}
�"t�%SȂ?`��߰j�A�n�"���W�h�글lc����9��bxj ��V����sX�>dʴ�L����ص�W�D,s�W$Z 0t���|G$������GM�=�Ƀ�&�����26�t��H�f0�\���n�Řf�݅�o���R�&�����|[�s� ��C��:���;��.K���^���r�F�4�Y*��~�N����ܛ}	�:J>�����-�ř��GǇw.���ߓW��i��w�z�d�]��n:h7��U�@;DMv8i�	R �"͍W�J*l~_��ū�u� �2�n.0���C�c�t���~�{B%���k|B�,��-Kn:���΀�s���lK3�����ao�>di�9D#=i����⣬G��4"l�6TTD�ON�la�b	�3�#!W`}�N���O���J�����Vw����K?�@���Xܿ�
�yO�E��i�NP�m<���$��y�>]"BH��Lt����dT������a����L��U�WZ�c�@�ࣜ�d�Q΁G��t0Б �Z�S�P(��Hmz,y[�9����m�����%2�w%�r��Q��e2�G �"��{��z+A��@���uD����rw��qj91݃6G+���I��䦃���C#��}jG%�z�%�u�`d,D��ڬ�߅=|/N#� W(��X�1�%Ih^4qĪn�W�!�̖��`�e�j!���O��C�C"4�D ���feô,]m� ��px���r��\>Zv�ˈ?���&�5}��k]Ÿ����͟+��fx�7%���bQtR�啍��ĞČ��r����h�Q�Dvd�}_
w(��H�H������x+�����VGa��Zy������p����SYV��.2s1�q._�#�^��6J�u���*�R��h�AQMG��\�<
7�sI㡯P��?�jW<��D:ކ�#�%��5�nS�!UqRm��� h3ߖ-?���ei��#.%MF[�z��@�T�A" 5=��,a.=�O�;��iVoXV�J"hx�@��xgtC"����ǉ�����e�V��}c��� l�f>��sL�n�
?�c�mb�����gB�%/I��wC%�$�\V��5]�ŵ_UL�w�k*���LN�j-�9h�}g��sY^ ��	s#Ԛ�t��l=�ǩ���k�j[6˝��0:�hp��vi;R���0�����_����B��7[O���{?duC1�������x^bgo����`��w�]�+<��*��^�
a#���B����]L3@l�;�0���Q��#	 켜���_p�MCi��[[��P�UJ-��z>o��c� _�iE���rJBA����ф���"�����y�p�?��~��bw�ul:0kQ�TL9����ƽ�7(��#�c '���T˵;�C��c_v�虗��Ɲ�N�g�X%a�|��5z(.�q�^�8�m�64eg�$�|6	��uqk�4$ƹ䢽j�
�Q1#�iL9Y�C8�)C�\�6�)��lTd�ab��AЛ6K�DmZ�3#l�<�e�s6��l�c^�UJ�(�\H�{Y��;�i83	�C=p=\����@{��{�?��q�s?z��*g���aW�Ʌ=�,�7G�'H�1�"�HsHJm�/["3�<�sj[�ٳdp����Ƽ���T�M�6GN{���)�C*��!ہ�Jl�κ�ɀ�7��� C�f��t���'�h"�]C_���$���c���?���ɾp@�vĔ|��&݃���g�s,n�(�u��U�>Q��M���ߌqKd�0dӶ�H��3ES��.e:�t�E��{����=�Y�&6�F̡��GA��Ο��z�[�͔��q�{Y���W�Q�6�Y����R�B�#N���7�ܞ���KW� ��({%JnF쥪6k��zy5%�x$+���:��g�x�ǹna���@���%�*`��,z�d�߱|.�,n��x�I�P�01 ���aU�֍#��$dX>OF��E��й	�i{�a'y��=L���� N����'v9�U�M.��f��u��H��}�z���!��q���5$ʿ�7&U��\j� �p 3�-��-U-�F��0Bn�L�8���A���9}�(�) � iv}���c5<�p�A��c��q��LH�o�îk����>���Ԋ�ʮ�҉A�*�<�b
����Td�\`��e�CZ��_j��ɬ��O��[��D��`�]�n�Z�P�N�{��Є]�F��x��e�6�4pp��dA⛄�4���{��f'��]˯�ሁ9_��|�D��-��\=3�B�|�e�T��(�Q'�� �5�r����1Vh���~객����)���!>3�'RG`�H����%R�W~��RE� f�I�ވC<�RZ?�~�W��*��H�t�;��u�Q�G���
�3c�	��?�-��}$'�M:�����0��۝PF��v�
�J�T��C�K�}Z�3z3������L���Dn�r�Y��D-L���Cݯ��ڟ�v��5=BH�v�ݬ�K����8ϜBh�~�"!����b�G,��R4��>�-�MT�!�n6���iQ<�b���:d�͕�����.t(���Y����!Ʉa7R�㌓��-�j���`�(;6H�rv	x=�4�X��y��<j8J����p1�'�4hVz�#�m.?0���b~1��L��\��.�K�6��BWҳ��vم���F���m`�F��p���"��A�M�h���< ��T$�t6�}��wQЌ�sD�М:�nH�����v�<q���;��?�@fZ�%#���֐P F��H�c7/�)ާ����޳y߰�W�O�<�O���ܰ�z�I�)ʻi�����P���1�4��E���2�$��_����m�~�&�?�*~�4�X0�a#+��Pt�otg��H��s��[ze-���yf+
�w�������G�t�h�ު���W$L�>܆T'�22�Y&�?A������&1�(�h�o�za��o���.-^tvKq����N]m�t��1�*�:9���j]Z���i�ֱ����{�@���F�҃�G�8Sr}�~��z����x�d���@���]}������O�;��D�� eb���b�(������M+n�[��ݺO�`9���Y�N�~��j9=d�[�Bt`��́���S�-��f��8BӒ�È!�_��X`�9�8���[�DYƺ�<����&A���6)	����J�ؽ��`����0��.Y6�����¾�ÍK8�4���LtP�Õ5j�k.����h��G�{����i��U�u i�P�S�fl�&lI0�ON�\��c��}�Сo���ڊ�g/�/�P�G�G�[����	�?]m�"�t��{�~��"����v�cU��@T���z��y� h�p￀ {�}�Q�L��e�@��u 6�
[sA�����mt�;���PX���&E���n���
����uA2���
���|u���p�c�����S�,>���һ��p�Xy/R�/�ƚ���䂇��J�#n�k㤄=���\�W��]���q�Fˉ��u�]%�ا� ��p���>�2���K����1�[��ֹ�q<P˷��yF�lj����;�'�4��OH�~K�TU�a��T��k�Wq�2���EZϺ�z��	��{3A���(�H��Y�V"F]}�<d���|h�."kzݾ�������P����c̓@0��||B�v�6�	$��~ӵ���pQ���j���(q?m��v��a0���0�����`�&}8G��͢�mVP�����5V�rf�'�a|�wĜ���/���u�j̪�W���.|�Vf?���	WJ!m��ʤ��Е���+%6���T��R`�O�yg�.1d!ѨI�Y��*9����]f?(ܵ�O�c[>E!(����f��jSk�r�`\��>#�|>u��I��(��Jb
ؕ��Vڈg�4I�!�iҮ��.�n�n#I"6�~�d��Y��}���Y'��h܀�6���q�nr�g�m���J�W��>���&R#���֐B(�ĸ�rH_� �z���$�r*쟴�Oi�B�!r8�9#��=��[��X��d�mU���2q�˦���1\}�Ed���)P�7%Tw���JU&���@�Q.d�3Hv��{p�e�a��`"��z��I�e�\KQH� Į-H����o7�~Y�C�i�@�����W�����k
Z8(����^�A��S�
=�S	�<_P��W�Zy�,�~/��*�r��JHF��3�be���kѻފ`yH�gUF����sS@�"~G�M-Z�3nF�M�q�^�������]�:t��u,�Tp\cM�.:��d�\E�Pi%�aL�c�ݒ.��Er�56szFwVK���P�>G$ꏮ����a�Ly�n�,��yH��
��X{V����`�*�������:�L�}�cmo�aF�i����@y�o�W�q�I�6�p��/����֜4��൯<L)q�$M��+b�+0&7��~�p�,�7+�&�p�7|୊����`ʠM%� վ�q�T�?���1	� ����G��Yd�q� N]�,�U�,�3�j5b����=4�\��;��:�f� �J�ݏ�f
2[�Y,�:<�� d��c��'{l-z��'�a�|���/&T���0O���ݼ�J,�7��t.��;�0
z?\��RY�Ŵ�:�޸Jy(�ݸwm��fAZSQCƶp�4����MDqj8Z>�(�n�8R�Ҧ�3ǟ�����^xG��.���(�X��"�\���[�f��6J�������´g%�I��j��{w��C�v�2>70�M�a���?�M��.�Lb8��	�f"؈o�6�]V��c�r1N�cP�9R����L�����!�����D��@��*�ԡ�[s	���p��Y�q�|(���C�UĆ�֧�D3u&j�N��V)������	�(�D��*��W��pVJ	;#�\I1������j ��p�{�z��5�`mz�|����(�J)W~���<�)dh��o�A��:�~�V�"��u��s����b�Ӣ�R���Ma�&,k���%U��͢�d����~���X���i�w��Jw�����HBF�=}���NsK��e��Y\2�G���V����|TYDN
�A2�8`ɴ�"ߠs{)���"�:�@]��G��6-�V�S�WE�8�ޘeNidí�ݔ��,;M�j�Y1�=�� �PL�W��xw�	ً]�3B��{r��0X��\�:Z��CL�=�\2�디��\��6+�� �ȡ�8zCH<]���%+,\F�4iP��8V�?z��`!|��K�=$�|��rf�z�#K�fK=��g[]n�8V%	��U�y��)��]I~T����o>��K
t˪�Z֞ s\��\�3�Oh�o���b�
j���:�j������N�����5���=�6qZ���a � @�\y ���P�0Z!`�e��C�6qg��T.uW���=�HpZ���z�QU"��q�I�O��ea��H�i�C��%����E`.v7T�*��r q�X�e�y���{�֎��M_�7Y�Dj�vz���8j���g��\JJ@ɖ�1�'�+mI����_Y̪�n� ��c�B�F�1Q�G������mW�x%XWPd�h��?����s1z��z�t��O�oK�[~���{5'F=���Ƣo�ZM۷l���X�_^Oa����#ԪU>1����.3q��(_�(}�?��$*�T�T��^pj��}�vG_@���o�ۅ�b�q5��SE�K�r��j���7���k9�z��x�#��q82��WLJ���C��6��mp�g�V�a0L�d�J����c\��_j�5��Gw+M8�2d���m'��)"Vx��_ޡ�AQ�Ҩ:�_�aEnT��E�w���A�����cUiS�Ҩ��6��Ex-�� ړ(���J�l0�:���?��^�1:�Q>�^���k�셿<��:IF7��`�uP�+l3��y�%�l���+��l��@���O$��S�V�2}.��P��Y׬�N�'M�~�8�H�J�u^�L:o��bQ�n ��ڀ{���&���Me[���#Zm��3��Il&'S\@x�騂�#�gao����A]�H��fL�I�N���&K.p^�R.K�O�x]�\�g�E�1��`�����>��t��Y4��7nʡd���-��%'�iK��T��d�wχd323ǫ�k7UdtQ�o#F�G[��&'bc��y`t�8&�$��?ɍ|̂՘�a��LFF
��Ӻ�`ϙe��v��B63Wa�k܆��n��������2VOz�jidt�P��(8U���{56Q'�m~�MU�\��
���b(Ly���t�?wM�n�q��u���C#�{����;�yLBϫ�����a�e'ٯ�v��oy�M�i��iq)��@�{Z��o"Mº���b�(� �zҳ**��.�r|�VٴJ|�^l g��	������m|�L>�S�E3��x�;!�)m7�@����!*U��7X�T�PL7%��.��!�>�T{$7�+(����tG_.B5N��c�Ңoݓ)	 ��2Whr����u���it�R3��)"�����@S}�Ԕ��X��N����#T }�<�=�8��㷨��o^K�C��^oz�۞�?�^W�lQ��B��>��˿�̙�2h�}�$$fJ�O�����;�T���e	�4�RՊyl8�|��]��AZ+�����I�V���M8�gO�u�]Q�jHb"�����J��W�m�K�6��*�E=�ot!/[�a�/C�*m�s�H�Zt��e�J`�G�42x���+�#���8�xD�3�;"F�/ %7�!���)��_j�cjξ��.ZY��}�.�Y��/Y7Xr�F�{b+���eÈ��0��|o���y�bn��8%��eNd�g��	9l�;��i�¡9rؑȍnI�oR�����gެ�IL�uĒ��5�����/�.�br���!�����-�E�^u�;p.N ����#L�I��(�7�"AeVu�yF��� O6�]���l��)�5m��i����F|~�R�23-�C9|����il�oUg�̖�᪦z��m��;�"������H�����oS7 ~���u���[����_

zk^��n����]��R�h3��v�Y����j@Yd�t����<"_ӥN{����tJ�����QĩZa�yx�<�>�~� ��I6���2	���M"�=D��ڟ��3��x#z}��PY4!����å�����z�����f����p3�'�`��~������3����ҵ�=ݫ�=��o�w�:=80����A
�N�����UJt��-Qy�Y�,��k�En��j�9��׼��4o^¾����cͤ�,�{W�(���F�c�W�6�*���_�fx��U�ǂ�7��t9�K���f�cرCz��!ݼA8���i�D�����7W�\�K��7x_�+���B�lW���\����P~�-��q��0
v�.�KS(�RR�������98mn�.����ݗ�`� SD���t�S�|�0٤��T��ٞ���Uۯ�����8��M��l^�&[�I���HYwqp9���0R戯�͍�L'j��}�������Q; DiS����nx��EڈH_��OI�-J���D�q2ٛl����*�sX�X��Y��=���6s!#�[~��U*�����B�nT���x���W�I�kh���i��!��4s&�,�ѯV\�/�si6�`�\����sP�8�بH�ӓ�Y>,�Ѽ�Z��a�a[��).��ZJ�p<�����)Y[��I��?��~��}n>��w����70aX4v��)���h���V��H���x�Î]9lwB/�2��1�<�lӦ���V�[���;������4�gV4e;+�X��k�b���+�5���Upѥ�q��F�&ia}�����u#/�����H����^2����͙3�}�ҥ:���p�%ٵ5f��K
���/�B�D�~ې�����p6h�A�sV��.0�t+k��Y�9�d_i�����X3>(I@-"�[��Uy�����ZT.��"�y��4�Ԛ���Q**,9I�r��d�H�|pҥh�m�o[�+e_�q�ԅ������#��U��#�F[ ����{l��/�K\�J]1���6O�P��k�^�����k����<i�mqc�/Ay�M�\p��bޟ���s�!���嬻�����}�Wj�=��%q�\����[f��Rn��~mȿ17�s�:�(�����î�^HIy��Fe�t�Ҥ�p������A�w���R�<�BW���i����AH5'��w%}TBQ,��-��~E�s̤Vc����T�$"�z��@���H�Ɏ |�����ab_�r1M�s
�k^���. �3���� ��������i�]��a�~�5�M8_Qؽ��DK�o3zD�>_��%�1��F�,0�FlP�O7W7X���j�XCEB�{~sJ�dx�[~D�ғ��"�������ha��T��������ފ�S�p��}wjw�ot�v����R�T �9��f�!r9	�~��a���)��r�F|X�=dmz�=���bN��t������}�8dܝ��9|�W�ו�LSTT��[%����`N+��qg����`�;��:����W+�M���i\BT�zlu�赻L��l(!�-��d|�/JB�}�e�Kc�(��<�r<~���#����������}j�䒞Ub��%#�Z4x��!�|��H�3�b�`��}�S(W �D/��fUj�p�:�T�vb������x�6�sn�� 8O��d���Q@':��D���&�gK�����>ࣛ���Ӭ�sٟQ�Rئ}m�]4$��B��� �n:��"�gm�'��w^�,L�f)a�.���^ų�shgBk����q�K�i�!"��I-��BJ^)�RJ��E!λ�ǌ���>����**}r�����@)����]���9@$����{�����dR*c�}���>����`RECKЙ˒��ř���תxDRm1��7�L�u�?u���S%����Ú�PEs�K^fiE�P�RgK�h� L��l z�礢C��Zh�.+�g������Zʍ@�@�0Z/WbN7�X3�V�ڿdt|�oL��=;���ᢺ����2M��=��(��"�\lv]�3���v>�tYNYT��]T�gz6�\�,��1���Ƅ2�1F<����f���d4���\��t��;Z�f�����;�������/u�9��\
о��D����h��\�/���,5�� 0�U%��(▏�������픳I̩> �J�?���;�� ��pW�/Th�3��9��La��w���R��h^�"m��_Ӄ��)ݠ�<�J���Uy�)Uo�	�U�h� ��$e:8�z��0���E 
*�2��&]�m �vʮ�!K��,<����N�s�H�߂���йW��[�N�3�|76Ң��z3NN��_��E�u�"&F)5�b�s)�@9�F�9���b4;5�o4PS�.Zp���ؽ��I�Ui��+Bn�+9gQ�0�w�Ce��Lr���b2���8�9&�~j�ni���;q}����kUʥ��z���E~s�}��C�R �/0�q�'��W�v�_�=JK�m�.���;pg/P�i��!iDh .��$+M��f����!/��&�6=�3i
�MG�Q�[�K�%�t��fvz�#��m�3	]"ف<��io��a-˃4����5���T5���!6��F~o��;���R����},w���j���f�_��pu�h���e��ֿ�sH~څǾ'�����E�0Ц^��r:�byONI�M-��9gN���qV/���+C��[���_�MfC�ܝʲ�eN�����D�{�&�yO��dn����dl�${��OX#������vd�l�����A#�{��0�����u8ҋ�3������2�2����}��������ݽsט�t*r?��0Їy��C�!ۢ��qF��Ɖ�NY�B�ɲ0j�ֆ}�W�ٓi��Ċ�H�5iq,5f�1�<.!�w�� X���Qy7#��|2�Bɨ�{�{�"�� �-�WF��܂<�sN$!��#s¾�n�yo�j'���&���>�3��|S��m�#�W�H5r�b�	������f�-�Ȯt�^��)��f�8[_>-�Hj eL0�>*��B��BCƤ�OjH1���r���c��yʳ��K�Iv�gڅ��q�F��ৢ��zC7����+�T�>����Mb'q�ֿ�Cqǲ���^�2c���.��!�a����ʺ���k��v�300��nh~���0Z���HB% qO�J�T͵��y���C��޴�NZ��c�/�"�Me�RX>LdCc��AR>;'��ͽ�.�ǉ�)�=�t��aĵ���%���6w�K� �z�E�i�׹�+H�>�.h���b6�՗�"0~l�1ڋ�K�Q�!�ۡ+�@�T�H?�S��fwҟ���έ%Av���1��5�-qy��,�5�5M@��o�:&J0L��)f�|�'HQ4Uu1/��0�D�8���L_!�=�>��ؖ��)�k�`?"�?�BO�yܳ�P7�)�^hE2:�z�����=��A�v��"��:K5B��x?ձ�Hb_�#b�-h���/3.+�?����o�aQw)�_15�l��^�Z���EW���H�ڑ�nݍW�}��|b����[ԙ�å 2��lCiv"6U�vC�jr��KI�_F���ie��Ə��\f�R s�3����&H�]��ϴ��h�)y��n�1_H���/�d��k;�l�W�|u��/���xW7￱����W�������ƀ����|���s7R��I�	���X��Z �_[�L#��oZ�ץ��Xs����[?��� W,���uM�A4R��g�j�S_�xw��3�إ����M��J�������apUj�\����yP��]�j,2�j����;���[f�3%���u/I��O�&-�B�;��oJ����Kȩ|XHY�1��L<x �Mv�ZlN����!�~�lk;N��;��ׯf(���[�A=�6�������|X��D����M-��Ͷ�'��Q�i�hzO�C�fA��<]݃��"-�f�}x�^�B�R� L��'�9ڔ��_�zU�Z9��1��RG8�d[6�%�K�0 5Ƒ\�l3@�p�x)��V)����hQ��h�c�Ї3dʄ1�Z8��dĻ�����(���D0'�0�Ps���f�'�q��n~�{8W˪KH牟#?&ol5Sb��\�2�M�����,r��tJ�e��Z'���Qx7b4}"[�,-O)z<�d�F���rI
�9�+m�P׫oZˠ�3�y�~Y(G>�����h�G7����=iPz���D�U��zV�3�٣e@�?�=�����3��<p�8��Ϡ�[o�_��#~�g�I>_����]ͲA?��f�3Q�m=H
X�y�@�B��"�믌m��$���������x$c5fk�b��}��q�p!�����S
�z��������N�����z��TP�}8ٰ;�b�np.,�ş˳���/@�E�]�%e��x}g/�wA�Q|5�`K%@��.fF���
{`,.ac��sƵ���K]��rE夎�����U�_���(��ǔ7) ?ڢCE��	v(߈0$��m�U��P����y+�����H����
���$�=Y��A�w_Y?�g�*���M��!����iN��q3g�o>�/}�qC7�!ĶE9��X$:f<j���@4e����hߞkD"�uM�?J�`ȯ���pK.m�T�&{��{�tz�)�<�|B.)}Va"�����
���F��J|R�p���΃��^��1�����KS[�׻A"��F�]��qL��w�����H�lL �Uw�t�BR�����Gbڵ�
��C�*'Z���e��=|��U!$Ɨ~�ƺ8u���K��:����+�� ���`���z�o���-Å���Њ�]��š�m�Y�T)�:���`T?�����U�\�3�?�A��#t8p����$$ܭ8z,��C�֙��v��� �N�ӥ#�Е��DT�$B��*��
����� ]D8���yXM9ONZSѦ��;�IN����|�z��L..��q	ANɣ�H����+�I/�l�a����;��;�_��_��8���H��G�a��}������Jް�W�{Q��hI��T;Q$� �u��&����: ��;���x�_yGG5��p�\�3�"a�x������R>�_8\�4���ӟ��E����"�Gs�҆��JUT#7x
DN)u�a@�f^Z�:�G����F|�ޝ{��^l�jQ1��R����A����Z��ȁ�yA������CH)���l�q"����>��zS��?���{8k��i�]Z�W�B*y��2���S���J�W{��0����6��� S�2�P^ ������㎹+�x�_����٧(�?�!YG-D�l��9Š]�ζ}@�kp!��/���	1 �\dzy)�t����	{�ǂ��%yE1;�f���>E�ޗ���!_�	<���ɥ�\ب�_̓��H-Tb��Gpd�-��$:p�"8�E�0R��0Z��Y)Д��l�3E!�R��y�yY��=ן��!;��D2�Ҿ~WCkc� 3����U��UV?"�vг1qtI�𨦋�����<iL�6�O��1���s�(ɴGV"��OX�y�2�i����q��^C�b���e��[���I+����u�ȅ�-���X�g�Τ,k��(55ml�U{�2.��s����x�+��Wh�D[h�J�±��l��	e����e�K]�{�i1�up���`Ioy�0��� �qXe}�/3�vҀ3�9���ymF2�̭~�wۍ/�$��$����6�$NRF��$��W:��WSxw//����T/��1��}쓑^�Ƥjh1r�צ�'x���F+��j�����OI�'���T�v��U����E���ŉѣp�.�����醘eT�á�w��d���h��?����w���y��"�r�R�������Z�D�Iu|�ܹ*-�W��$Ҍ}��<�^Tt��\�.�\2�%/b��������EP&ύ�3u���8��S�|1�X�e*�k	b8�Fq�u�@�e�m�7�L���Ts��ī�l?��8�� a5�I�"��Ie鬗>o�|�_(?]C����i�A6�����c�@a8V��L�=�h���@&����t�[b�k���HAlv[dbXV9e|x�:"T������]>�ڰA+��W�l�@-]T�
\'���Mߖ(��r�R	����^Tܒ����� ��[��T(X��N�O��?;T7�����ҷ*&��[�N#����%�䍖Z1�u�.>,sޓVk���Q�x�HA:_K�0����QLV���3����%芳99�[<��[���I��n2��J��9���~(*[��!�#�m~O��]r@�6�gemo�����r�^�=o�ӷ�R�ul���Y�|�h�G1��c���!� ��I�#N,ª ͌��1~�B2���f�rGF��~I�M�`E��~�m�!x3�VH_��.Ǐ�}�|�94�#�dT����'O�c�|2#e신<���W�˒�p�=��t@��\��r�n�Uc)���S�Ɲ-�do�������J�D�#����_8��H�5˻Oe�j�y)��mP%дe�Q,ϔ$���[�!��D:��4����)��[��>���U#����q<�S4]�Ǧ��C�'+,qc��3K�|�%T@d=�@��ȶJ���R��Nn����~k}��ThǕ�(��X2��X�'	��>�R�r�N�o�$�`�(j�P 7��U��oqo?\&RjI��9��=1�z�3(1�j�L�S1���r�f����'�BK�	����{���:ܝ�1Tq��	�T7��'�ߖL�XCCM3�7�����}�5�Lze�Ј��;.H"��%n �.qq����[�RR�l��n�Ќm1���O��p4W��:��}`&���'{������u(z�� �� �܉[�^3f_p����n�щӵD4Z��6��F�D%O��{�E����-��#-e�@O\f�o�ʄ�|�h͒ok�N_Fc��#�s}s.B� iG�&�	��ُRmP���×�.���x>,mܹ��ű�m��1��9�u,�^�=N�������Ѱ����0�ǘ2�Zp�0oP�D����8ѥJ�#by\;#�~&�x���N�G��^���V�l�V�e9�^VX�����X��G�Ɣ���hOǀ�a�<���цub�8�_#�z�@H��{�A�(q�q�ܜH�P�7��V��$I�Qկ�
Y^򼶗W������C�<���'�1Q�_K���	�!�c����� p.jV�D��A�����I�b��2r�M��#@��E�IԿ%,e���BÁk�@�C�k���B�L"�Ǹ�H�!�u�����)��n�"�챍O��d2�%�4�~���Ȭ0���Pس� 
�F3�@@@a����rw�E��Y���k8���U�Mi�B�C�\5+㒅��Bf����@\��.���[.�-��3#�$�Ҽza����U�OK�CG��r*_:a�އx�ү<ȥ
��*�U�Z\`o�Ν��|�Ԩ�ߧ�7ɏ���-�¨�����CAb��'a������0h+5h����iv��f��SU�A����<�RP|Z۹6w��s|�&P�W>t��P���+��Wy楜�bڨ���g���Rg� �r�qdJ��i�:�^]A�ߓ�g�3�@�_��i�#�y�u5cs4�2�0�Gq��BU����<�g4Sr�L���Z����<;9��K�Iv(���w ���1ɡ�b�\���<����x��CPY�ZW5fW[���ꜱ��"@ӱ�t����&:�O���tfF��+̾�*�$ıs��
�<�N���?����4�[�B�Ycl.\Z۔u����mJ�.���a|����Ru,~c��>E��R3KI��2��O{�R���)�j^���e!�w�O��F� ��W�u~����ۜ�vb�]�.�����%�*�o�dܻ�O/<c��!�VDr�U����#t����v���y ?�x��V\Շ?S��5`w�q��LJ�&��9�QiQ�%z�>`A���@4k%�9c������t����4��V���`��x�?S���J@�O�þm�%�L{,=�Ǎal�1�Q��~�������_�H��K Vs=9`Jx�+�PK�yf�>w�m^~i$��M$�h�K�	 �H��`5 ^�7R�ɢ2r�u�Nؿ�E �tN�q56<Q8R	i{Id�7l�>H'ow^�x���J��j]�*%���I���9'�0�\0�W�fڌ~V�˘۵r.�P�Z[��2P��^�5*�L�sv�B?�.�2��˥$�9�]c�/X�dw�[\;�����ZD*1�߃�Mc!٠��9�N��|`��0��%
.q� ���a[��q�o��ȝ���a�mTP�⥗��9�|W�)���{]J���q����[���b��zE���_ŠK�Efw��>�Ƨ� ���"����ȓ�h��<XX��?-SU�?`+��C����a�<X�L��lgk�2�O�S�f�s,�4����͞�>CQ�wYp0���0���}
�#YՊ�DaZ}����&��H�[웏���`���`F���t�mC�H�/$M���^<H�f��=���1` d�Y�����uI|�(���\(�n��갶zT:_sg����҉�4������M]�6&g�ݠ��R:��әsōxDH�P�nN-�A܍D�t�Ӳ�Eui?j��/ʘ7��:vRG��p��[0�T��5��$���O���H,>�#�����շ\^�tiY�ţq,1r��KR)4����S��J��O�]��Q�	�l$�w>��4�`�RR<�_�#p!-h%i9+�p0��=�P�ARW��/�,'���!Iw����JFcS�Y��)�k�t�51ȕ�a<��%�ݣ��tO廩�V�Q�K'=t4GU�= ��������
��$\����Esr�T�|�&�����Ɗ� !(�<����{TKT1J�X:��K��;�9���Tu8[&� ׇ�c��$6")�J�WǮ�9u#��.Š�'=�#z�SE�S"��\�����N^ٜ���o��/j"�cK7tϻ3N]����pc{��y�\�PQ@�x�j�ВX�K��d�bb>��IMP�گ.\V��3�|���O�:ی�|��\�jX���}C&q;�*n�[]�X5c�!̛P�]�g9����~c3��.�x8>[IKQ�ӊ����d����)p܌^[�#/L�fb�[���7��D@d��3�Zشʥ��JE�V��$x���q��� ߚ�t�r)@H��$�	u�R��}м�B�%����A���:����f�3$�;a? 7<<V<K��Zt"%�˧�A$���& ���;j���V�ĴoҼ5M�"sx��F��1A��|3����B�����f��\�2�"#�}�ÆZԄZZkƎ�x�pi)�[����X��פ�Ah!߆��(<�p��Ո�Sb�6�?m�p�n��|�q��$�O�ր�?�FS�������6����x�k8�P���6z�5��,��⧠���s�٤_X%TU�k��sJ4*{�'�t�}' (�B	Me���ޡz�]z�$֭HJr�O���AƵ���h&n3SV��$O�Q�ә�|��!E�u�4�s�#�o��|-�΍X�(�9��m�Sr��W/���i9M�:&F�"�P����ב��Y7*Uݰ:������2����#w�?kꐹ���5�6|�G
�%a���薈�z���ܰ�A�݋x8�~f�|�*�f�k����zҥhgF�.]�j��݆����}3rw�
��;җ��~E��y�N���,ӆ@�n3���\�K���lyy��Rg�(}Ņ�X��h	N��W\����ROx���@uS��s��J�ִm��O�G��F���@y�HJn�m���p_v�B�g�s�Z�W����e�wq��'+Iq�)�+-p��K���>~��|�>���[�l�����$����8��T<X�?�:L�y��ñ��]pK���ńL�5��L�d09H�1��w������|�H���#�K�RhA9���b�8�e)�'k0��c�/���ZF<��z�ִ�l�PU��^�!TJ��DD�~�2�Dv���Ηt�O�Dl Hl�"�J}O�Sy�UX\�0ν���C"�F���*e��^si�����1Zl����``�4u� �շ3�g�1}���#��Y��*Ct��G�>�C_]�#�?�k:���`\�ؔ����9�1�ҳ����f���ę��fm1��o�Clɟp\}yfj�QѮ���m�y�$����x��� Y�3 ���Zg�Ŵ��c��!;�w��I]��7�69y��=��U)�c���ZZ���^!��n��W\S6Q�y�Z�{)<MDZ^A���o���3 �t� ܷb������i��,�֋��x�7E�U�����c��W�̀k�0UO�P��U���q�@?]b���._ ���U�Mg����kRi���Ueߺ�E�M���1s�v�����ʉ
�$��0b�Wj���O1�L�%)�a �)Pt�Q���5�C�����!�I����(�����.g�F�Ġǹ~��`���҄��j�������pX�05/[��,�e�/�PY�*�[�ib]��nJJ��ɉ!n��x�XF0C-����{F�ay�/���v�	�ȱ�f�x�~>��~�"��I�9N?~�]q��k�E�G�>`�m�%�t(sM�a����s-56:��#+���X�
�����VPp��L�}BF՚L�/��&��m������Q��I�^Kq���w�~	d�p�o�i\s*�i�1/�N��o�h��t����)՗֥�Cd�<ǒYr�Κ�o���#9Y�6���f�R�j��iu׋,�6�o���*�C`���c�%�Gת� `aO!Q���3-�#Q���S_zj-���G�N�	U[��-O|h?�;Z�GhY��+=�7Ɏ~Qx�7�OαA6�r���?�i➵��5
���n4�Va�FGK7�9Xn��^!�*N��Z�>���۝��,U+U) Ѷ�)rP�����v����_F��P�X�R���}2E�GB�I�KT�Q��V��
M�4��*�/T��?����.�!����RMx�e鷟�џS	@P����ېp�䕒g�U
oɰZ�ϒ��M;5s��V�Z@;�L��$AƏ[~2O�ҏȢu�`�Ә�}Z���01�B��	/?X��f��0�Ϋ�0�={y�34��2�C�ʺ���OU�a�C�[9%��XN�+7��Zi��I̝�L���/ ז�ZCj"� �u��F��*drn�UdQ�&�P�"��$m�� >Е݅!#r\����Zq�n�5uK-��.�]Em	L}����+h`\���;VC.1���q�B��䡆H�TE;<f�����q �xJֶ�>\��
r+l��oD�l��(�K�6^g	R�V�����6&;���r��\�}u�$&wKb|M��P)�ػ�	ZP��S��p'F���n�5c�u�&��c
����z��Ñ��~�\4��㗕���s1R���َ0�睑���!/R��T��Dz{l�j�Egg��1ed��g����C���_�E�0��%��/ץ7�����%��!I����Q�C���&,RD�?��$�p!f&y>�����Nb��|/9�I;n*�=��S��,Y���K�f�5A�eH`��5�^%�>��r���oբ�զ}�Oc�o���j��}�$�O]�*��0l��}�X���$	G:�
bz�E�e����s�k�Bx<��m�7���tp:0^�`�rި�"�+��X���1'����V����!R�Oi��$�zНR���a�oQT)�h�*�V�ϮPjy�oM��^�x���Nhǥ
�2��'�G����f��ƹ��Z �XJ���T��	h��y�;�F���Q1`�d�;od���z�w�>b�lf�_w�-��OH�}�KDmy�7��pH���T��Z˼�̳O����� �B���t�G7 !<\J��uZzf�N�Xf�G���/g�3"��g�!wv�^v� ��/��~u�T�I����&8�����v#��m���\����d_�W �诣�Ԥu��$<>�̵������AQ9��̠e�wP|Q*���/�brA��,A�&�E��L�� p������\eL���Z<�ܿ~�>�6�Q�t�F��U�*�`�)��?���O��CPԢ=q�ۃ���;��8�U�1�f{���y�����K�7K���!�L��A�)�Sd���dt0Ad��:V������w����"��MZM��Z�{j������R�����{}���:@h� ��~𹧀z�˅kD�,�U���}D�ц|D�8��HqӋ���MƱ�V|x��qxL�����@��v��U��?�qi�#�~��T
bee��n����N�h�Y�%�IЂ����MJ?1����[��S���Ӧ�������;�dv{8`�&R���3��
d	:a�F����2����~W�'i�%��Wˏ�]�]iȟ��x8����x�_� �@��q'�!\����DwK#����I��55��Þ�f���y��M��]�`D���]>7�'��� ������ݳ�< �³���w�1\1\b5P��6��p���U?�ڇ�L�x[�A�. �$A�M>R��F��u���y7�"o]�c���Dv�v�
�[��w�y�]�5� l;ȻM�:��Ǳ����/�̲�� P�9a�?%J'G�s�>ɧ�kT�tn=F�$	�Z�&Aq}��ւB�b���	��'ITS̿W!�Iw6�Ih�r�zbP���]���:vk�;/m���NT����*,�!������E��"3đX��T%;bQ���3+G����(/��K*��4;��~1�����T�ć���� g��4(��B�":�15�k�e4�����FE�E"#;M�m����l�:�V���F��~�����b <"�7�h	a�ȷ�'��$FTWQ	��O`Z�FK����Z�����C�վG�/���@ܑv��,�	)G����!���G#��!`,\����i>�=��Sȃ:8�����՞�J� ND��z���㴲��k�u��RB��Nk+�=vy�i�}o!՛�^?�ze�q&/�󂔱�l>��K�Sc�C����	����K^�B�~6ɤ߂��`4�в5W�p�`Ym�SA⓮��j���w ��N�m)�7y˙2�.�����eQ$({��U�n1�)_��n˒���o�n��9�#'ɝa{��$Z�"*�������
H���	|��!_B�7��i�RPжOo2|L-ߋ| �V�����1!��1���<W�r�!DT��l������Z��ښUfË	�t,	��Z�&���ɛ�RaS5�k�)G��ċ�����D�X�_&Vb�ĐU-�w�陕*��_1������p��S�3O��'b#������˧'���e�)���h!�)�Q�kQ'�*��P��#�kE�X���{d~��D�ċ�*���߰n�k!��4���0�d3��޾\|c���_�.V\p�$ɣ"�������j� ��46"l:��i䟾8����)I��%fG]_��X���ܿBpy���c���ߣI�+7���M�qV�/����GLN����܍�:8#�Al͙z��/H����G�q��T3IaZ��#�,���|���Eʆ��Nn����?��Boh�1(gf�G�D2n:�u�w�־�w`���:��҆_i1�g,mb��¡�8%����<�TIIā��s�U�Z�:��3��O"ږ�tS��
�Փj�c	/�����O��.�<#��e �� BBnN
5/c�R;�L��~��j��D�^�����;�}�s�*��4�E:3�6_aGc�ikY�=:�5W7��`����=͢���n~d��d����+j����jMToד�+�J�Ԇ1|��L�dAl�SghK(��dhK1����ɼn�S=��?:�F��^��(*���y���e���m����;�����_���&Fτ�f�~\�"��X��e�D[�#�n�'�#U!eg�<jĴ\֖�I}�T���\@�͚�+"o6?������$�"�/�ɘ8��s6����]�`�Ωmۨk�k�j�3`m�0Oz��}HX>'���}��9���fڧ����9{��M},�s��JS5�Y�#bX/ԽF���̖O�!�)�'3��A�b�l݆��z�#�]`l���$�Y�Mү�Dq�ή�Wx�v[�U����6�a�"�7GN���(��T̋y��XUl����aq�G��NDE��
�H �aE[ AP�+�v�6�ܗ��_������E;RB-R7�3 ��'��h��9����88k��_��;{8,!����~~[
Tav����'�42�}o2xȨ1�bԁ}��r*������x���Zh� �?!JH���&
9��3'�5U�"%�2�_�<����z&�NT� �����;� G�-�{�LF�$��F�T��ȕ)7���O�ڛ�%'U�:�M�9_5U��\ %�>�)^�]E<f]�?���H��P���:��6�9���DX����d)2'�li��^']^�e�r3tw;�#+e�2<���M�h��T��d�[_�:u'9����;�_���fx�("I�/&	|GR���������M��=���n?67JT�Y��F���&�r�u'a0�!����&U�k!ː��R�Z���X'<uEg{	؛|W�e�c:����^<7IB���~���w�QG�o�2������$ƻ�����$�1��� _�0R�d"�x�(���L��T�Y�EI:%YLM�8�]c`�$����d4���9tQ��85��k�zXv9r�h0H�
�)�A�Cc��o����Ҕ	o�!^5�9>W�j�>�n��q�ڜ0m�Ǌ?o��Ui����b� eh���Tx;`~����e{��pq]X��<	E����kT���e�C��r�w�A��,+���E���^���!�p&9�ԋ�p��d�z7ѱ�r�A���i�#�ur^����BJ���XP����J0qbt)p���A��uN��>0\L�)���)��py��U���K%xs֙��#��Č���C	�L媅'�	\]#�����	�r�3���׺��0�A��+��d��o�\C-����,�U��R��2~ΏI��͕�)�to.���y�g�S�F������R�U�td?��Ǣ��r�wY���K��~��d�0�9�ihJ�P����U��M˃.~P䤾��4��rUbX�5M6��]�%4�@�ފ�(�R�v-����7�꯴~���j��Rd����Iԧ�-j#G8�
���=XQXX7�c�^(���K�r6�-�e�A�N	+�I�mR[�A�S��p%�>kƕ�４��`ȱӞ�����a]	�6ƴ�rD��@�A���|�@�h	�J���͟�U�xTC�=�4��{D3U����J+bH�^3T�#�#���:���"{�� my/PR�ʥ����ia���[�u�"��с6���\���d�Y�ǘ�o�-���^�o��;JY�%x���S]�8ɡ���;�����a��d3�j���1m���=��{�G����1���õ�S�>�:�&�[�O�U7��A�#L|)��_s�.C�a��D���i�Xh�)����9Cw/�h�S�������y�ǐ_�@Ie�>�嘱�*?K�0H�(G�X�]��M"�Te]���٣l{hAs֋�c�;�����gN��8R�E��J���rN����bd��^���5��X��>(S�@��Ա� ����$]�PN���	G� �,��3��XD>�d7��n~ť%�N�?����㧩�o9��s����3�W���B�� ��hT�"���W�����rhz�$�/8e�`}�V����%�u|�3�~U38�� D������f�\�F|� �5�5�}|�f���������Y#����|.d�VJ!d��u�4�UYh�ON�=J�FO)�+ųG�L�R��G�\ӄq�$/�
�ڑH���z���Z������c�?� �qS"EU��+e؜�&�>Yc�&"�m�;�yP*h;�����u��X���  ��8ūJg�^�HD<�G����-�ۘʊ��MSK�Y��0�9�� ������]�p2��S+��ѯ��N�XmB��X�����o["r�Đ�u�F��=���8?XdtL?"�ҍ�Wb�F
�_?�{�k=J;a[QG�+�����|����q}����9�L]B�> 0u�v��L��y���>�J���э��@0m4U����.o�2M%~=Zo��n{�lB"$S�:K�i��mN����!&���Dk81v9�܁]���Ξ��I�6�e�[M)�ls��
J�D����'�ԧ�
4d����LO+���?`Մ|�$N�c�<�����@��h��st�Ǚ��AC�.v5�چ�ǽ�>.-�@d�P�f���#�Z/9�������*Y���8߽E��]8��<|Ȣ>��qL$8Q���(E1��1��1^} ��
?b7��4�i��lJ�f�Ye�z�s �wP���Й#.�l6 \���v�՟��q�jn�^�3��'�A�l�^#�VvM �kU:5E�-A�2��Iş{(��D�̦�F�n�A��z�	�˞�?���|LEh�卛-y�����5;!-b�&�DX���8NN ����Τ�~ �d����k�)j��$qm��z�Aņ�V���V��-��_J(�.�E>�#�� l�V�Ѡ ���O���Yg$���c�-5�\�����,ZG��n�IU@TW���6ӭ^���X���N!��4���'��v�g��*��]�E�,��f�ʓ-��am�*,��{֓�@BW���⩹�%�d;����w[M.9��X��'��v=�k�u|�[�19.ߒ+�V�:y�� D��8�}a��y��x֒��#(�̵���:���(�n���*sg����mf�ܺu?{�*Bj�;G�n3���e��4,%��$2�d6-���J���͌���z���K�����'(��W/SLW]�z�5�㲅T}��U����ۡ��&l�$�8$x��t�6&�b.�~qq��q�8v��:h#t�J�쩭k��r��~�@:ã��H��n�ʌ���D(��qI8��u�ј���m\�!l�Nܺi�L��ސ=uKf���Ax�Z�NVk���k@	S�~�--��Iy�= ��ʆ�ŹqF�d({5�k[��H_�Y�d�u���tc��H'|m7�BU�ѫg:y�<tVO�\(�	t-�F�m>��/��T:��&(�o{U6yM�CUP���{��M�Q�s!1�:pN�H�r�Hى��}s��ܺ'��5��U�Z�5�i?]S�+��$�E6z��|�:Ò��d#�,�	�"d�MA�MѶJ���C�r��Y�Ќ�N`��E����c�o�����)q�?K���ߝǈ�[?0U���bb`��0w6u�B� I�=�K ��r`;�丌���E��wu���J�j��4�3s��u�) ��,s�2}���$l����Tt�4>�5�Ǣ!����Z�/�jbB���L�EMY����.�U{�v�YOו~��0����8X&4�!}�m�!~��T��)F�����ɡ��.3ň;|���{aUR]W���`��0ȣ?�Dץ�m��GS�5䫹Y�ih�킨��7a�j��>IS��i���*;eGF�Z �ژox�1j�,��˷���Gp�`�����U@~|�1}Z@�J���r��?!�xʔ<̚���1�W��0F���b�"��u���Q񐜚W�����4Z��[�J�� �4Ə�TX_�vdX���m�[f� q ���a�h,�}~K�1�Tc�++���P��Ƿ[�`,�8<�B�K��ۭ�:�<�F�+ï��[(��}}G�[Y��aфRk�����=���\��}y�����d���U��1�^m
��?�%��	�<�l�F8e�n���@��<T����v�R�2���G���Bc���Q����X���Ԍ�jʛ��CN#��$�5����f��
o�����0�-\���l�%�Ƅ�b��4U�_o�D�,��0�i���5��a���>�� JZ��� � �#�<-7��PE���up�uyXu|V̗�%KK��M5:Exߨ^�,$�2	�S�4�\�5,�g##�;���i4�Kk8�� Q���>V�eN��]=���1�~��s[������?	��v.(���M5��*xSk��g�5���Y�(�����#��+�7"��CIW-��(�x��M+��!���L���Rq
��ʽ����\A(�X�,��U��ל�dz�p\�Y�I������$}�in�~�~*<�Y��U0���JF#���3��}�ѢGBE�ν����Q0w�>��^���=�AD��җ>܋�M�� #~Nc��-����-�" +9r0���G���9�����8�|���9�"Z(��ӄ�J�7Y� �3��߈h��]�� ȳ�OwsM��V̌WYu��>#��A�0\�h�js��/W5�@$���܎6DF9����vax !���O�e.����<). V�6g,]��yN�J�W�a�*� d#���olYC� ��LL0��o3���ؽ(s�Aڝ��K�6��s�fJ<W��N�#�/�Z��[��ZsE�+����:���AA ����K![p��)٠ժ>�;�Eb8��E�*�;�|=��&6t�3���m�ɥU;�:�����R���Ē�J����7Ͽ��g�맄�2�"e��a��$����ӭ���iQ���~�7'�gD{����m{,?m�B-5> �oAeFvT�k�<���|QyQ�Q�*�G���R��+�:��ՉmqR���Ҫ"�tuw��3)�>� ���v)�C�T��ȅ� n���wW��5���1�!��P� ?:|�@�,��:İ?�c�Y�2���(CnrN�)�a�{�h�@��l��A(�#�&ۆzR�S��3����Ӂb���D��ԇ?4e��#���+K��WE� n�%̌A�e��F�q��h��-1��o~D�َ�'M7+j�!F`�)W:c%��&s��%�C@,Z{�s���� q�lP�a�����u�x�� Q"!O�p��,�ἥ�%O�,}�Պ~����`O���a��Q�\�&�9*���~���V�rS����?�fWS�E���ۍ9&5��׾!����\hRp�a-���Җ��ZK3n��1x��YK��o%^���7ڱ�2����@�x�o ��F�d�Z{���,�Ү������}�I�lA�Q�"�r����v`��0�����Az@�A�n+��7��F����	sJm�`"�'���;��&�7�1?�j;Y��ÿ�Ɣ�7E�
:����X�hVpZr��|%V-uY���Iy�V}g��\� �ʳ�X�	>����"��nv����"JԲ��PF	����[�0s���`�H�Ga�U�yr�k�!��>�!�U�V�}\F,Tܥ0y�A�g����2��k��a�ɴ���2�@4�@��Νꍅ2L���_7�1�������"�W����4h��C���ءp\c����Eן���M�Y�he���d�Ԫs�ڦ�����K�n	7V�L�� ȞB�OI`��|S���8�I�_iY�-9�`���Vt�5��F*������dɰK�c��t|�е��|5;dJ�C��RH��'#�٧�(L�h�?�a�����f5�$�X�_oh��ݡ�=���A���H)1's�L��T��#��K������uQ�*�p�T*���-���V�`��r�D�hj`��f���5�US���H��p��藜���~�����+�����Ѹ͝,��������*��e�%}[�)�� ����A�%���1ǐ<��o��}w��3s��E�F��a���
b{��{��m)�\���b��}f�j�Zd�"���Wu	[���Z��[�p{2� b*p6e0��,ɞ�uWOddY����\Pq&�W6>�r��"��J�"3����B-�Έ8\)[��b�n�B�
S��,y���-�7:�������O!��l����E��w2c�)��Z�]��Gg��5EP�zi)b�H1ml��b=E�^1����]z۴�]2�Jkd2�(�v� UfC�Fd����8�G�xB2��&Å3i��Lu��[Q�SS��6����cϿ-*-��h|�}:�4x���,t�C�  �:"�)��C>���[DCɢ��w[ӄϬ+E}�O��
�8���h� ��ёK�bD#�
	����E���{�{<���#3�+��z�����M��re˥%U��t�	P@Y�d�����TQ�Ď����
��K�G�8��9`ƻ�_��b(fi�A�=�]t=�L!������h'O<��Z���6�k��^(���smI�ƒ~�VLD��{�h؝���@�X=~'�G'�� �l�g5HǮ@�t;22�����Q�rt����B��^^4�ϼF�6�""����JS���汀����݌��'������ԉ���m �l�!d�]Й�)ڵ`&.�4u���x��C��>�=�P��\����PM�Z<ϷyY���2SV��������W��A���d��}�&�PtK߈{~.B�*O<.����R� &4�D�%�rXͤ�@�\~�Q�S�p��pa����r�bp�.G�'��k��z� 9�����J�]~�E}�(���P�Ox�Z/rk�`d���]�TxgY���2.���<��gP������P��o�����EU�[<�@|gm*��ͯ������:�e���'[��.�;/�Z\���/ `<q�,��juhw����Lz�<}�l�@u���8<y��&ɨ!�{^��X�Y�Fi4[MQ�����~�y��*p��"�����̹��W���hL��'��A���	I�����kn��3��[��]�OY�dM��X���f:�!`�w83F��B����ty�|��x�b������X �IF���9�����m�{��ߏ��k�TF�Mڣ����F{ɪ9(s�E~�i�[���^=k�)Db�h�{�J��U Z [_Bv��%�s	[�#7���6;���zE[��H�-&��y��@{iA�>xKO�9L���4 �1昈٥$��9Y�K�@�k��׫(���ޏ4�v���wv0��#S�P���I������	����{��6�����Y���0Դ��Կ��>�Ҧ)V�r���֢�dnT��_���s�HD�x�R�^�����.��&�f`�ۦ03�ce��>��\"��2�a��ll��A]��SUj�\�͒�_�Q�8�K�c���p��t6�� ��_��"n�y�V�^�����o݊�(�6��(�VMo�<H��]85�(w��0v��mI��o,��7e���̯^�-l?��5�(�����
m�
)���)M��*����-��*(�p$��1�Ǭ�R���g*��%�����O��tDx��(��%6 wwC������g�1Ƈ�� ��Q>)��J��3deW`9ʽ��ۅ~'�t�x���d��IZ�܂����H5%�YX�C�����\n$#�C	�)��q2��n���ưal����89Y<��n�S�g�#��
Y������V��ѩd�T0������~�m��j�E�
e�_�F{��YSh���E����<�wr�'�T�v,��U�%�I0;�d%G�Q�n����F�>d�@�� ��Z�l«/lA�gr��B�x���`P7�:KƋ��F����IB�*�VwG���	�o������G�V_oxd��/�J���E�dQfy,_�Ӭ$��M5�4|��H�Q+(��߆S"s!#�P�f�`�����j?|��ƹ<���\�HV�X5�ey�|�?$Μ���z�?�w��0�̡�;+����)�"ʧ�>�9�~Mo�� >�uUHHQ8HD�~nYp�t�o*?�_���Zǎ�g���ɓ\�i����B�0&\7pVmTFh�I�����T���S�Tv,����aC0��|��B\�L#h.��� ���SE�ӱȀ� w+�=@���0�W� ���������y�<��T��՚�,��wޖ����/Y�S�T`ud�;�X8U�5�b���4���]�A7Y'\R�P��h1�˄ �gc5���й7��6`���ҏ{D����Ïw�1C^4En:�5 5�-/Wi�����d��`¦|�WVr��pa!��Zr��QRў�y�DĴ��C���I؈Z
��K����B�XE3_�.%I�n\y��������Zb}�����h�7;
�6>VnИ�'�\��Z�i�fbT���� ��ƕ�al�XQ�Rք먥3j^�NT1\���UT�t-����Q�I'ۈؾ��������`��gR}�x�ofP6}\�]��|�]�4�
@T�.��^4���w�Y֛�l�@���5vMf��TM�����G�ʹV�"�B~H�j�/y
չ~�_%�uÄD�l���R��$����ŞA�����簢��T�@f�����D��f�|_@�&|S�����Y^\
�pw����E�ڣ��~����S5�*����f}��Hl���~rPTWKunB�/� ��,���vH���� � r?!���M�����=�{���s�d���!$����u�e(1S���[=ܞB�G�XV��!��ĳ�y�DX!����C�P�h���ù��64�H�J�ߧ����1����G�Z��b���[�NC������65FS�t�����s��F:AP�-���Q�nR�I1+�[��Y�:�^�7��'��dUԎ�%�9}[�g�R�I@Yqa��h6U`�\��r%�E0�k���t�䇗`��%��yM�@,H��U���D�t3��L<R+�0��)e��c���8n����\n�~$������	m4�tz	��g_%j�oB�����������D��e��F��f��U��5���=�&	�����Xz�DX�lH--�ό������A^#�!�w̶�?��-F2"�J�"Js�Ͱ������DrM�q0����P+z"��J��S��pX���$WvՈ\��?@����AJ�Z��-�~qو���^%gB��&�F�t���L[9I< �\�D�^.�UyD���L��Wk�bs}\5�\�\gxҡ�9�+g�;�vGm�T�Y�jN�4jo���Q�_�Se�������n)��E��]�U�݁m���K<��G�E1�ȉ"l�E�&ROˆ��
�!�LG��Z�$��|��0�� g�N�%�ƙ��JJx4ne���b��Xa}p�c-���Q��$]rZ�F����e�q �S$�`^���ݧ�K �/ʽ������33�����	�T��o?P��=�T{�-!��� �a�"+}5�x�Bc�̯�8��OQ�zÏ���J�8�,.��@�u0D���])q[��	��Q�����\�Stx�-l�h�B��R�q�[6IW*�vk��2M�+�{�xEg:]+�q�D4u��7&�Jf2;x}�/}�����[�m��@{������
I��k�����(�MoGl�c�C��b��ҷ=��<c�²}����]q�mƾ�T��L��t�p	��m��F�ܥ�vl��$,�L�2�x-@7����
QU��2<0J�#��D��>7�נ�݆Q�c�n�ODQ�A٬�T7�6�a9�Ԇ@��>%�W�����BN/Յ����XMo���D�X��审�glB;ٝ+c~�],C�mԞ�+ z]y+�����$PB�ӱ���0I�p}*ܨ$֛nλ	�3��1{��	�Ed�Q�Δ)X��S��;�6�9����gC��Gh�N��^���@vv���G���dPd�qOU�W��ޝ�(���0 G���%y�ğ��vB���x�2��Pi���t����a�u��􈵄-H�Q��������)|�jP�g�ĄZ��	�"�%'����$�YB�I�X���4`M�s��ל&١ΏX+��PR�`��	��>�SrlB4�4>��x#�)����d�Y�;��+����Cn��69���7�'�:W�05�6�µ�8�N�QFqĒkdE,�,D�#��)�1��.g�P~�Q��Tp�o����2�4�'�<K�)ZC�ӧTq�{���!B�TQrm��r�Ą�]o��0�E�_�J�<v� �P�9��|��6]YWK[��@J�i9�J��~m�7�0�P1Z�k�G�+��ր1��	���N���R����0���@��C���l$�w�r�Fx��姣4}�sLm,��H1'�J�V{��������N�vu�a��uW�)Ƀqt�]�*��y�m�����23W_�8�Z��p�D���p[)A�W��l{�²-}�'::B�k���U���#�/�*��~�Q빑t�)��[��H'yKI���%��&?��ć(���|9Bb�������k�'��W��Ј�`+_�U�d۰�8P�!�h>�����E�P;����!��rsWhXO� 3P�Ji��y.��kb�G�LX�R��S�q5�~���֊�V,l<����Ťh��#n����gH��\z�1S8+]N������(�Xy�#Kw]g��T-�V��]BI��t�ҹ���ʌ [��#���ks�2 �n
A����İ�3�� �б�D
[d|��bZ��&�Y�$�#�w졬��W/�^�T��N��<J�Ԑ{�G���C���P�`�я�!�g&��b�l0*ף$C2X��e�;r������*��evt�0�6U_�j/S���P>���y�/b71�YT1���؞�r;�1=o�:��ܗ�b�v����_c����5�צ�J:0�2��6Y�~<�����1�7�B8��C��C�MNr���XL9)�6���2��Ω��/N ��V%5eB�T,��0�~>��2C�s��گ���f�G�W9G�9۷��c~�xpl��?5�7#���[��^"*Ny.ȷ=����1�2��e�S��1�K�{��� ę&����E�G�9��ÆUy����H�����bWyV�֤���Vy�*��]bі$0֯����mh����y�=_ʚif��ȥ�1�[)��F���&� �~�2�z��rIfOYaI��PqD:e�X�0��k����&����q�L$s��m�5E�N:{J�Ƞyz�\�����R1�l�b��ȩ ��A�����g4cYK/��./?�kj1�@W���z�z)N��u1�ܣd:��6���Q �49H�܌HPh��i�0}�'�/p����j����4�UZ�pw�zH�F��c�	b���\��%� f�bSb�o	��⟴�d#��R��z[e�\�K+�]؈�GmHUE逻?�ljH�����g�m�x���F�r��} �t��$#��ph^N��#O���L{'y�<��V��B!�_�� ��'u��#��˺t��3/]$z�[�e��o8�!��Cʮ�X�]���G��"�5_{��	�L!?e�rz.����v�i��*DO��8��!V�Nb�4��f���]�3C�4�	J2���k�(ÓUf�Ѥ������}�F�6SZ��<�QJ�U�����5_���oC�8*Rx"��#���Kr���i���m�$��Y'{�]���'JNUӨ���E�"I��!j ��Ȼm�F�$pvJG���MjQ��Y�Re�|ה�bj`�g y�o핯�A�/ ����� �a3N��u�.I~5:+`�O�C�.��-�30�w�h�M�"��U����$ݛ�f7!.�*� �P"�6���74m�Q�2%���CM�n$8�j>�{����L���2���i1�F�r��ո�pa����-]�톐�QB&���!f!��inˮ�^�yV;���Y�+�j�Sߖ-=�m�m ��5P�@�<�SeTt�����X�q���]����تO=�(�r�$�W��d\}Ve�0#E ��f�z�Gb붊�����J�;�=�)��)�J��fP��[h������%�j�孨$��!��b�8x4�(�M��3q�l2�U���;�c�?~Ռ�x��`T����v�(EwI��j���i��Ѡ�U��bEY�Y�M�N.���,�W=f�w]RA�� ��j5B��%�`g�J�N�uM����(A�u�d�^2;�K��� ��s��c��)4P��� :x�{Dq�m��b�8�S�`��K�&�J.�s뀪-�cw�3��ˎ�:�GA�ܨI��b��)5�6^���*n��;�_�\U� h�S[:�G%��BHe�Ô+Pt|W���/O$ԃ��#\u5
��";�S;/�lm��9	;�/���b�C�]m�WE������ם�G���.~�Fd$�gX�۠�OA������:�m�<>�R�6�j-LB$��n�7I!��{:L�v<K)M��]L	9
���e�[�=�f@�j�2*�91U	���
g܃bF/���򆞓��b[��갱'�jR%�2qV4i���Qָ��n�0���/��{����&� -t�d���YKG g3�B�`WFu|;��C�Q:�H ���v�A��4'���>ɑ�~C,̌��9�/QFuf,y�����j_@\�>jx�-;6?����J���� IW4��$P`	�{���W������ou�G���R(J[@��ef�����<dD`Y��Ra�iUB��7���v"����v��~8���B��>�{1���S��,�T\�7��[M*$?�ޫs�z��6/��6��*p�IO�6A��@�M.�T�P¾*-3S6e�)"��&��ZծO峈���_�#�OnZ:���%k��ݸ!Ʉ�t���>�������U�0�y��d�+#A� ޥ��J�<^.Ad{�k)\�[	Ri-MN�# �,1"4�y`R�d8���Ƅa�*'n��	�%�]g )������e��",����[��bj'��ݭ��V!9	 ���C���>��8i��%�Ԭ��&�{F����W�Fl|�l�mT�
g���/�A�%?��
��r�'��#q����U/L�H]J�Wl
/n�5��l�δ=�G�Ԟc���8K�ߩ>̛�_ק�h!Q��B�����4���1U�Eś��8wH�UF�!u�]y�o�#�S��v�)[]�!�����U���<)������@Xs�Pm�k���I	���A`=Y\�c�q�k�)�&�bLP	U#��/�0,}h����4���$+�#Z�'UsYo�'�_VY���s��]F�� �<�M�i#be�{�YE].E�l�+�>��6�P�g!���~��7��l#و����&{� dY�@�Ǟ'HU�sL�,�Y�ͪշ�Q3^ܭ6�;>�>�2��
���Ղ�/��5��a�sM��$�U���wí��"d��|���/i���RE#�� ��ў�||��65�٬���mC�ƞn6W؅��uM߆����a�M���\PMB/�ͿW���F�a%��M��M�,h�uc��DC� H�hU�Qz�z�R��uwBtY��.���OZ��sh�W	��Cy�<c�<U���O�Z3u���+�dGJ���t�խɚ0ͨ�'w�R^ە���F�A.\��R�~�4�|һa�HE�@�9��\� �f�'���4��"�pg��k(��h�f|�+�m�i�d��ґ�>,(<`}<�=��]�"N��ƬQ��ne�~�7\��><N��;ᒚ���6����~�A^��gJG�RL�E;&y���0�#�b��s�2aQ.G{�уrb�����Ow�AY����X�>�+�f�8N�:�ŉ�/��Ba��^^v
�&��}��'ሥbv��� 7������[��`�{�b5�^V�x�t�~� �bπ3��NY�����~�%������Hz/��$Y��Rh*p-��s.��M���wf�U�@�B�o�%�^~wU�����J�����$�x�qfv��8���`D����F�Q���^x ʾ��|�2���Tz��02]鱋_iu6;).��7��%+S�B�l�7�4�� <������z`�[��A��L���Z���sܹ|��7&�N�>��tó���I?0%В%�5:�"��Xy��&}=ce�W��s���8m����Ѳ.Rx�wp���[]Ğ�;g8=vҸ��	��9^evY�KZT L�[E�e��,��m��C����]k��2�i-����ӯ�,\�Q�$�J���r�5	%���HeZF.��,Q�쐪d�鈛�R��} �R�cʙ�ǘ���p�:+v�g�ZuE���A�g+d�V.�dp���P7Q1mn?�}���?Pf��n����&8={#e�1���}�,*eRDRbv#�O�3����>ӱ�	j�(��EI���=���Z[N[[>���i�ќ^]Ʒ�X�t�x6F�����W�V{��qTӸN�.���� p�<�QI�1H�sb���5�[ͣ���k�.=�8 ��oeM�J�j5���&t в�~��M�+��\���z�W[�H��"E&^t�t�e�+�(ۊ��v�'��/ئ��OO,ψIJ��eѕ9n�Q)?vŀ�a��Xӗ>�̊�bꚳ$�Zc�"W1��}�k^�	��0S4���'���D�/���>e�6���_�����"b�ըѦ
���l���P�}�h���~aq�����{x��_����ߕ��8��A��a��R� h�~&��H���)��3�e6-��.����(y��y2_>�W�\x�e�ֈ%�a㹓��R�Pa�/o�N��_�zԜ��u��_�XwwʼO�wq�M��O[���z��tg �7#!���
��+�^3 ���Q���"�2�f-���u�5Ѩ��9�#ݼUv�)ZWK���r}�#&$�9}���Wz���y�D��a��p������+3���N1��~�}��M- f�`F���r����ʻ�o.���m�'�"�0f~q%e�5Z���>��`�M��������|�*�/1�T�^�	T]��v�"5��~�|���X��i��K֐�4��	���Zy�6�ROǤ�g�������^L�[<j�k� <�Ǣ��%!S(/F�mX.r�'������<4�:ϼO�F����m��5?�C�7���%�{��)\ɩ�\@x��Y�2�w�Äg:B%�t����-J��;�jcgI�a�}톛���k#nʁ���\%"	�YC0���ȆyL�W7좈$w�`��[�6o��,1G�i���c��7��t"텛X�O�Uo���<|�f������)�ӫ|:��J�����~������������o��^<�w�3�����o�C	Q�~ l��ܛ���7�ۃư|�;�^�y���]�CkN���e�����Y��5]�b5��b�n^��4ڢ�"���
b����Z_T%,
/E7��~��Z s�
o�>�Iok���LA��qG59��Vs�NT��5�C�l��a$n%�����Ig��/MNLr���$ �%�j^7��Ǭ׸Q��	+�s<|�>���n�����%�UP�q�0�����$v��Cc����~�'Ֆ>[6�JE*�hY#�5��D82_����`V�B^C��f_���"w�M[`fKW��vT�l�W�h�</�i��pi����|О�T?zh�>��d���&[�t�p�Xtt��9P��u5�����5�s^��h�!��x��C�$�#�5���3�Ǐ���<p��έ5<\����m��,��>��4,��e�����S`�V��d�A)�͇����ʈ�A׵�M��&���2�ٻ-r�1Έ�0 4���j�9'�1k�u ��e��s�I�Ⓩ2�>��{@�-�K�� �Y��򬔓i�~�р70��8�w�TK=���R�CQ���5�O�A�ޯ��&�����&�!��+�9*$��λ�H��n���,�@����Yj ��vq*紮��QqO�j��TVP'!J�^��@�DJ�Uq�QOB��Bg6�W!]���l��O::C�0���nm�~%�{�a]Zkr.HǴ��w����{��ث�d�ܗ�IV'�����q�$�GJp�C��>]�M_\��Go���0F&{Z����4,@��8OPӺ9��įP��"�HՉ��+o�.!�ɬ^��$/���l���C-R�3�N��X���L���<��xY]��m�5Ҥ��� �U����k>�iJd�������9~)B�7�j�S1��(Md��N�H�f��ůDΏ�iG]�9( ӒZb�ۺj����ɔt2z^s�M-\ �@������Z��8��Ϲ�vE���Ԟ�4�K��w��V��Y�2��2	�$�n�Vf �摫Rx�)��.C��%�[O�f�d-�O�B�]���!Pe]K�n��X�i5��q���CU����Z�w0@�g�^fa��F`���lw�7J��-�G֮�����8���]4�[0ݱr�e�"��'�h�m]��Q����\	���|�&>;�4��a&�N��]���RAPPL1Ţ���	��*\��7�ơ�3�J��;����ה�}��5��	P��Sn�~Zu
ө6C�1���@���E&>*��5$6O���ņ^Z(Κ���R��܎N���F}���qlW����~2ȑ��Cw���Җ���85 X�=���?At�@�+�.��f��&��#_�P>�}�¢�e��$أe����,ްF�La�Ee��L2����7�"WTkoW|�B@+FvWj�o�`6��zf��*�d�2Wʧ�@d���vR+���+��������/}��%�3m�����q��!� �	F*ws�$s!��2w� �3Y��i�^T�͂����<�aP�������嬞�<g�h�p��{��M����G\��kk:�;z�-@�Os��C[��c���t/>�[-�G�]��8�D�7�e����rM�R���ӗMҌ��>�n]��B,4�O�Dtw�k4ש��Ar��8_B�U�ǀ,V��o�j�T��%�*`����J�q�Qel%D8��m��C�R)�L8��֖�%�X�t������b���f�x�)�T8�=Qq�f���.
��b�A��bRg��E��������?;q̥����=�d���@���2�cБ�w����5Ŋ�r��=�ǫ>�{n� IF�Sޒ��*i�8�Rڈ�V�X EH��4����^�]�2%�-�zn�(�t���-&*E�JkCS�L���J�-��9L���lk��G�U-�.z�SH*�h�*T���)��qD�
w{��N�rk����ȱh��no��+h�."^� F�FX���R�H��|(4���2QSZύ��u�t[0 TT:��<&a�
�:
�0��:�.	���XR)+J�;��	��
B���m4����+t�0MW>/��<G�ԯ_!R���k�~Is	�o�9�c�!}V���y��5 � ���;o�;	3KM4}_�}�9L�OO���i���aO�|� $~k��R	�Z�%��[�w�p�|�6ƻ-��br���7q�?�Z������$̮����.HO��Gۘ�\�����܊�B��N���N'�6D Y�|��=��ym�8�����UBH����ˋ�(��K��Q�Ш,�$H�<ǡ�^���62����*`��\e� %�����B���yD�6�/T�q�w�=Vk�8n��T 9�t�	�ű��J�F�7 HJ��'E^<u��7�ԍ��Td$	�GO��B;�&a��H<Q���L�`��˻5��x!��3^�vf�EqS1��m��a�O^��sR�&\[};qb�0V�:�{J���h6�����YJ�!��3>x/M2����"�Eد�9'�����3�v���"7��G�/=�p�+,�X��x	٦��<ϱI�t�P7rW�a܊eX��!))^�6��X��l'R�~���-R�4Y�慆/`�X ��Y��Dm�;|z��Ҡ??H$&dR/雼�(��hjChTn��Y�S'��w�%^�B��g�66�Q�ˊ�(�9!6�Z���bn��7<�c��By��B��E�a��	�K1������Ϭ��Ȳ�,�J^�*��4ӧ�uњQ�kVM[c-}�[���Y�ǲ�O͈��ƪ��D���H@���9��c�˹c��d�J��^��`��*�����rű1�b�j5屾�\��hʀ6�'�&�+�R_[���R#�
�v�i�f�`h�1��Md�U�󼅬�!n!c��"�㞆��zA��4�%�1�ɠ� �Q֭I*�_c\�2Ψ�zDr���p�4M�&�d�����[n�у�y��;
n�m��#,�nU�*U��o��X6SH{���n�?�ay�,�.|8�wi��=%-��g�	O��8�� MYҞ��O�~c}vptC���SӃb�"!#w��^�n`�i�K	��?Lϒ>����P.�QJ[���H���9����(p�q$3���_/�Q]��'<3�@G��A1�'�7��d+k�\�Y0C��K�Ѵ����x�S@�/˂���z�7��9�SX�S`�nF���Sv�B�S�!�4S���g��+�u���l�-�saJ������LP�#�Y�Ӷ��qV�ע���	h�)�j~��$�U��p���d�����[Z�iE��x�?)�l�x��ɔ�����l�F��bb"�Ư��I��2�c�Ϝ���|�iD�<�O�|���؛����F/.����I�ƣ�hB:-�)��
��ig���Yf����'�Ě�����i�
	�� ����Up`M�a`�_]5O5���u�-��l?8}!}���s�9�B#v�Ձ�e�ʪ�u�]r��9'?V?r�Q ����w���"~���|�
T"�S��GG��S�E�X,bag:"�M�<���d	����D`ł��-��ٞ�d�N$b�4]�J���#�Nrˌw���a�US�'�q�пj�|bI�y�n��=i�p�x���(��zvju���>��e�r�h���-�^�9 B�
AS��yw��m�ᢙ����o���rk��V� ��K�5�Ʈ�v���� ��.�K=�������,�BRe�e
1T����=�(*k�1�{�zOl1ϧ!c!-���:�U'�]��R�;IP�.b+#�[9�y�e��Q`2��0=�6�*�����8��!�CX����=�Ŕ��E
�h�_�:�_�۟���T����9@A��q'�m��RM��sJ�� ��P�4�<���ː�P��hj��?�	��r�v���*,���z5��4�8��"Ő&���s��ֺ�P_��x��D��Q�u��~���js݁�jM�*1��^sP�x�����97t�iw�����R�_���+�16f֜ �g���"UN���	E0S:�dQ�~s_�I6ר9MS	'�T��#�<��������������V�/��p��Q>?�h�-F��(�
Q�d��ײR�e&�*~���O �^9�Z_R�_�Y�m��k����Q�%�7�ͥ����� �iI#��[���M��N��1p�A(��u06e�S�.ܾ�+e�`S�����;�����-�j0�N�dE�@m�x$}V�#��r���ρg<�E}�؄#��H�ŉvL��ȵ����^ y<��ȷ΢��%�{��ݩwu�r�3�?}��;]�V����ns�ا�~r�S�퇸VǨj@gä-��l��<a�a�׼
�>ؔ=��2))�w|��ܬ��[\c~�o4��0��n���RF�[4Hhs�
�'���ȇ���"�]:��0���QT#_[���T��m\..'I��]7ߣ���fMK2�f��irc�	2�����,�׎K��5��T����m띄P�E	�YC��p�Ӎ*���Eqx��g��[���0 �Ub!�!;���Z2��x`��&��:E(I��%iO�ۨ��l�&��I޿y�e���L�y����!q�,�|]��x?}��Wi�����Z� �6�R��0�����e�>��$��!���������w��K,����	��T��������O���Y��@�?Y�Um����~r����nP�+�����9��`��z��K��gF�95��c�6�h�^~���%�.���Xr�{�,נ.�qqt�ë�c��ɱ�u�膰_7�]�B�Uh�|�bz�Օ�.���e��IM ���R�n����p��[2��LG̑fG�6F��@�͛3t�END�|�h��\�h�����JdOF]u$�FQ��]����m���P�܂�C� ���	�kj�L�.�馊����B8V���kh&x�4\9C��;�rŏ`�����`J%>�g����3�&>*s�Y�r��)i�����{ן�7�
Q���[@Po�@� L�@��6>��F�о��M��-p��J4��)�����^�S�B�>��p��q��IU��WO�к\��<�45Ű` ޭ;i,�c� �dFi��/�E� Q�u���W��04?x��0�y����Dc��ۉ5���ȩ�a�Y�_����I���}��swV�y�K^PK���X�<�ȸ��?<��"�M{�q}S��2��ꋍ�џ�:�������}@(\����3�OR&|1ˤz�!će��Pn��Mqe��;��5'�9谻��9����X�y4r�|U0�Ѹ{�Q��D�Γ
��fbI���Ȓܿ2����9�&�w[�f�)�ݲ�.٫v�2����߫A��k
۾8�
&����q� �/S�2t�k�f]^'�#�U��qڈtf��8�ۖ��d�٩ny�y�H���`x� ��uj�R�f:3qz*�iM2�&X�"�v�"2ܛe�x=l�h�
R���ٌ��pM������UAq���&�S�¼�i��g.8�ƥԹ��!�y���}�nM��� �f2��l-�-������⹲K�7Zt����ޣψ"�}E��qو#T2%]0K�l��)5_���A3����q��>&����_�B=�֕[���\�=7n����E����Oa�n�w�Mj���¬n��@��[����Hy�2~�`�A���]�<��Z6�Ջeҵ������nWpZ�WW ?0�'�R�]GZыxz6.�pwt"��-8��u��;g�*S!��T�oH��ur׿�,"�گA1n��n�j��7�¼|TDz�#Ϗ�D�3��EO�\J�2R�a���e�����t  ���{x~�����3TO�!N1""�>@ݭ��J��
���pv[bsN#����?�g�|71����὘������E����>�O�~=mP���j����j�kq2I��`����(>	%v�EɵI�~G	�f�����'�D6�QgA��آ��mr
%X�j7z�	-�F%yƘ��$L`�AK%#�vuN��[�/	S�+'�����W𕛘�3�8̱<��5ϓb��&p��YͿR�N��C�n��d$�>����J�D)��L�J�z�����TV�ʌ5��!�H�"��|a�a樺[tb]��}���TJ���D[]�96�V�g�����\��LPi�G	Cy3�|y+���ޒY?6��LV��,s-@Ջ+���c�_�h��ЀX�؅gE�-y���9�zt��;���0%�	�������{@�?4���w\@
�A`�vb&�A�O]GR��m7w�!$̇��>��I��x��b�t�҇�7����y�{�z	>�2�q��]��9�;�����;�3O��)?��}��L@���t�{\l���u���l�7��̅�H�!�����ƃ{$#m�
��*&0 3Ҍ�/jY�V����7�ڍ.�¬@����2��\N�c9� �!y�G=¬�����8�g�I/��3M�����0��|�q˗J	P�>�P�?s����?��2��	ط�̕#������zs3�c�Z6v����D����W�	�'�
���NV�[n��5'�N1ݟm|:or���Z���5���ϩʦ�0TK��/��^�>��T�O��K(�A5�N����z�?��V��N���F)��^kg�'�F��t��4y����o��QN��KA�X�ؾd�y��Ң��>�aO�Y?C��y eխI�aO��NQml���Y��39�Oe
��<qE�9^�I�Z��<x7.T��A�3O��~�T���	��T��c�T��D^0�X���NtGY�Uf�[Y�E^ȄDOs�f���;*cs|-����(� �>Z��緘����Њ�o��g�e t�t�C*����T��J��Tρ�f&�nK�*n(<��6VhOq�z5�^�l�y������o��\���i���@�!��Q��i!�S&v�[����˅�m�u����[6�1�׳�y0>�c�y�ZU�WwXc� ��%eͤ�*Cz������1l�W���@������C�JV�?��HRbЙ�c��m�`{c������	V�\�Ĉ<
&>�A���qTL�]n��I7ux��y���c�ܑ�e�����1�ǘ����r\�K�T�F�w�85�{$e�Y���|�[¸'����������ˆx}��&N�w�h&��U�����ս��}{�w�I�&�C�Ͽ��Nl��<ۄCi���Ï4P[S���4t�z�,�	��8w�u9j �A�Q�m�1^'�/�qg��f��5�����e�u�ݯ�酪�*V'�i��K�w��B���Dὢm�-��ž��Y�$tW������/�7���<�e��;`xcH�4`��>rvT����^�a��x��K���E�J�B��"����*g\r�� c!t�|�6�l�	"�$��聯�]E������Ͳ  ٠8���Ð�S�m��NPr=�&�Z��1i���1#����؈���4e��i�y����}�B��J&�pjU}Е��T6��|�K��KZ��n�H�M.�֭�e(��$(stK��-�W��񨐣V\�����%TMBȰ��x�,��ǳ�0�������T�bO��ȮX�Ⱦ�֔�����K;P�j>��И����v�=A�1\a��;�ޟ��z�>#˾�2���"���uF�u����\j���	+Ux���\�,�]C^��Wy<���Ϝ.�g���/,F���K�=PUM��{���7�������50q���+z��l�ڦ�D:q��}���k�0�TC�^.`R�4"���.W�ͯ�����tN ��(u�����/th5-����O��#�r;5�4���q�'�1�&�"HV��1��:�XW;ޥ=��r���|�(7�/�� ���Bea���e�|C_�=��#���Ήw��t�����(������پ��x�1F��c@��@pp�������E���b3�n���� �0ݘ�zrH ���c��uK �SZN�B�O���*�{x<e��zg��>��l��t��D�](
����S�B|��P��.���������"/˶B6�e�D1@�~'�V{��:O3��Κ3�$w�Q'�:�ĩ\.�6��!o�J��W��l�R�F�?Uѓ���d�:0Qt�	�+1Q8OI��᭤l��8��[�7H����n�����E�\����~疥ɶ����r�K�d@�N@���9E{��P/yA��0�)��0�3�v"Np�φm�:N���A	��K��;7�8#��D��î�?���K-�uj����W��h�ePo���FQ0x�hm��'rF߂y��oҴ�;�o�@!"�]�?G��-pϾ�{��n�_� W��Lܢޱ����S��3��� �A��Q<�ʀ48���kU���a�-o���;��bZ�-�Y��"�R>^p�/v8	w0A}$�}
{�a�̪�l^��� �����[�ĭ��9Փ��o?5i3�t]�Fgݴ�(�����'ڜ:�Xҋ0�o����Pg�ـ-Uβ����&�����X���;h! ��3�.(��쨏�-�2�8��-H�_��A�Llr�DQ�
�=�l��C�K8z*���{h�ް	<�N�!�	�:'���i��M�PD*ޛ�f��Cg-�؆���;|"�9�jp�K/&.�ݐ}��ך���0����e>��Dg�3E�\^0�ޡ2_=�<�zh�6��N;\����p`/��QW��1Jq���Y�hpj�f��|ԟ�v�Z�L/9��YM��1��TzG5��I�9��1���RFHw��G�"��4��S��/z�xA��'�ģ�4�>�"BrE�}���r@� �/�rm�X\H2kI��[1W��|�r�(�;kD�6y�B���l���s}N���'ddp��AՊ�d}�g��s��9��òcVD���]���4H2�2:g«��9�>�� ���}����/����	�}��l"1��u�]�V��<}�>\	$�|����%�s󞕶a�(H�S��e��H�e[��N=ꪩ��%�8i3#�X�6�j�8-�	���ga��>��%�ftK�m�Q%���J$٩0V�/%�I���ƃ$ ���ѹI��e��d�I?>���h
�3�U2�?� ���bz(��g�C�o!m�w�c�	�7�Л(�ߺ㑻@��S�y��0#�?��Ph��Y�cMrZ���Q�?@��vJh{!�>�G��J��n*R�Ct6��E����"�� �_��\A��ỷ� }`v��;�PJ��a�	z����΀rH�BP�:��s��P��r%�ۂ�����tO��Ӏ��:������QR̸}�"L��]x�Ԏ]���w�X"~K�
ڭ}�}�UwA����g�=,�_;l��eH�JN�E�K�����;�h`��i�]fNt}oc@�o�S)�����d{5���Z����B#RhKt��$_7qR����:�kó��n��|���K.�x�2�N��3��ъ#�_�x*��|'��)���_1$dc����·½���:U��ʙ��P1n��J+)3����� �O��I�k�jy�3ό��LЙ��S��@��m<�H�C`]y�f���DE'�>��3��v�.̦uậ����)�(�^�c�t�?鰐8Tm9�9L��Ff�B��ض�-zo��8E¸�sT����z=s�3���ݭ���l����Xr��p<q4��o���_:��H�D��������U��K�.*��P�Z^��ϕXp�czi<"���$����_��M�_O�봹�n>`ح�V��T�{;!7;���Xv�c��ب|���_���T�8MC�\��!.B�L%Y�e����g(k��Q�G���D�@�G7P��o
`����4�6q��9 ��%-���!g?�8��|�W�N0��1ސ�kK�X���a*=�@�;�\�m��s�22|��+@jf���CI��%Y�|�D]%�SGj�e>�jY�r�I�F�x$�f`�S��_s�F-�4i[5L����ď,!��7�-k��;�ֵ���� !�h�֬�@Y&������p@�q�;E�;, ��5�ފiV��;�:3�#��G�M����&(f��6�"2��F�0��T�:�4(搫���.��:u�_�0k�';09T��0�;w�_JJ��Q�g�b2�oo������\"m�%hBt�r�ȧ�j���=�dmk��m���5�s�o�x��w_{\�RJ#n� ���@�Ҡ�pN$DD����� FK��^mFZ7���ɀm��p ��X���.���x/o�B* 6TA�c���ڰ��3��c	����:QAP�&�w�~6)�=�b�=4�"òf�M)�ȓ%��0W��j�l�:�_T��v���f66LB��I,�t�u��N1}-;iiiӊ�:-y[��y���� ��Y�2��g0-b˱X�k��xQ+��@�݉����.g�p}�D�CTF3K5�E��Cȥ���P$�A4����dWh�5b�������5�TXwFȽ	�ي��.U�π���Pa��z�L����MY��18�FL'����_b�h	����hU�I;��,��{�ǩ��x���y���l�>%�5�.�F�r��Z9C(��,��9�����kO�'?���mܕ�Ts��;�V$Z�Ժ5�96 �k�����IN|�CPC�|�|� �Tڸ�s�X����͋�K�t������W!��+�%�h.�
��B5�DW[ˑs�z8�_Q�fÃЁU^�S<���x)���9ג�APA���Uڦ;?�
j��f��˧� �G$�3�N���O
�;e���:`F���a\'��ɫ�[t��#� N�#q3a'�H��~e����?��O�Չ��9��L��L�io�!�@�T����bg�\�㑄�K8���x�$�§�5*�8q�,z�˫D$�e��ي�>D�T&*6s6�y[P���d
C�cU Y�*!U��d�q�3FE`��1�g�e�g��@e�%�=�A-�?=�")�=���4��������q+�Z��G.�"�vV���"�Xw����S��wP�y��̩&�f�x�}{�k"��*���\��}^�QZsV���d'j�s�:a^°6[G9])�f��,�[I����?upE�	�h��)`�rgq#����Fko[�JA]�E(���4�/�YeȖ�&�O>�K1���5��u�\��Տ���ˈN�"�ħtܪ��5�'ep^x���P=y��<����gw���pΐ�\{�'?7�����"�[���W/���?9ߜ����G��ǣ#����j�Q"0��y.�*��΅���$50��;U`�+�p�͜\$Hx�H¼����3����8�I�6~�"���N6�Z�x�f�_<��u�3��Lɳ�E7�/JS� �U%��,@������c��!}E�P����DI,"9G=��ɒ��H~c����
�%�﷧�i�}9��=���IY��z=ֶ�Ԏz��&�k9��d'(w�����t�"�Mv��� UN��r{�?B��G%6�@y�:��#ڑ&��bd�7N��hA���C�U�p|/n=�0�A���#2{�ű�i$�x�/g��X��;Ʋ׉u��8���5��I\����KW�g����(�eIa�OF4Y�����}�=��)��"�����J%�`b����@f5�6(���J���)<�c7��̣���ٳ���[�!Kg�`���&�������n��������M���>(I���h����L�{CU�u��}��VN�Q���Ͽ!�\��N����OM^ŭ/.-��.N\��_g�s�ǭO(���1� ���A�A8W��.)jP��7�muE��\�i΃��9����8E��h=����ۙ�|f?1ة�w%�0�����Y�v<�%��Ω�;�ĸ�I�yp~���ʏ>g�Ro�`��k�<�`�)�OG���Bg�	��B�%9b�ke��,eS@��ؘ�� JA�1�M댺̿�	�7M��h��܅��}�7%�\�0��=��x�Um��Q;���jݳAR �le�4S��hQ�\�Uv�W�#�¤���%���;:;����b�������� �C+Tg�XTX^��9��������U+�� ���0^=���\_~ޜ���.�R���i�_t-4�fP�׬����JkR
���ߠ*%� ��j�Z8bQ�y��{/���>k���XG�����q�O�c��W��XT L� �H�92+Z= ��(S[sr�̡�Ѹ�F�r�6����!�;rg����fc�6(�	�A��erp�!A�:�	�!U��_a0x8�ɮ���a$2�&��$cL�Ncz�Z��?P{ǹp���FN ��S:�����A�38�w��jԧ��z�� ��I"�J�u$���7��to͎��?�.K꼃D-��Ĩ(b_���R�ˌ�i�	ŭ_&�3-fH��p�H�(e��=���@�w>���?gR�:7�H���v��(��+��m��#4q'eL5����.:l9�b���.�t��v��$��x~��L��+<�O����,p�蚴��4��o�`j�DLk}}Q��:AZ�"�jil]�(yXd���V�i�)u��J�+���o#T�}g�}��ԣќRx��ҊxGO����NW���J��&�2�C>��Pf$l�?�_/��Ƕ]����C>[%.VVH�{(X,�+mC�M���ʪRe�^*�F[MD��}�jǴ�}p�OX@Q�����h?���U����[�c}�/[ѵ�JU�	]��y	p��޿�����px�U�f=��ɓ�ދ�O<���䃋�B�\���ƞ��S@A �}zBTD{���V?�~��M4��"i���C�r��F?�oΐ�r7����ߢ+(�0,�I�	�l�S�j2��°�g0H�)�r�(���!��,��r��mX+�o��8EDf_7YX�Sҫ��VWe�?X�)���;�{���c�XD�(E&�Lq >ut4��ŉ��)H������'��%��nل�6A���׽[���ד�W
�����>�_Y��.=r�����m�g	��ȅ���+��e�~����H����S� �$b���t(�Mt3TJ��ߪ�>]M����������U����q%:m��Ж�A=%��ϝ��Y	6H{`��3`6Knɫ��hVC������[Gq��k���#@���^�rd_�`8%
�w�#���K�����Y�۹+�6�F�&���o�;j�ˣ3|ȍ4^����9ʾ�ɌJt���-}�:�[����C���@S�_���=ӾD�&�}��h�y�1c%|b .�W��p����G�)&��Ujwq��Je�Nȹ[���ϝ��K ��3:0��G����wp>�,�z�d��8����A���d�ߙ H$��fz9p��9m6\�
�-�`^�瓍(�N
d�����!%����5���6VB7��F1��1s��h_��	m�u�[�:��ܦލͺn�v�������'M)���S����kS�yV����~�+��Dſ�ӫ�3맓fz�i��<TE
55������G+�l�Xֽ�^c���*�X���]st�k�<�x/�@G���U?�"C��Hԛ�mM!57��}}~�|ܱp�o�5����c�y
�u���X�ந�D�vP��Zl�(��d2�]c��(5 �+�Y0��q��	C�9���ך)�[�Q�8�9����&0 �ޞ���1W��ǽĚ���Bc h�l�ֈ/ʍ~����sڪ�h`����iȢg·!�c��׫EH+�t���85��������lZ�m�d���|*��ah��Å���S�����r�.P�9����F���ǐ�!3U?K�*���u{!+�_".<�Ù��]{'@>�����4q�ui,�3Y�"�,���ML�	5#>��9�	��{����.���~D�5�q��'��lUi�"�#�x��@����f3t{tr�W�.3�B`�4�<ދ+�2����y�=գ��h��%��-���s�c��
��HU��hB�#���an���
Ҷ$��7"��+u?�h�1��.����@���T�:�9�X�K"l0�3�)�f�n�-/e�':�9���̩�ec��c�	άCkp��~��x����X����mCD�v4�j���b��k�=�^�8���G ��߰���[uqU�t�,ҙS6� �U	6lBv}�𣔉�eM�ڜ�8kp���v����,�L�R�c�;��|m��i�"Q�8C#<y3h |����t��aɁ��{��Z#�=��_0]�=} 8��A���=P���|��>�RJ��f��l���c랲���֯�M�IN�-'���r�A�(a��Ɯ*�h,L��m+BD�q�/��+wDÊQ�K�*�U�� C��v���J��=5n����YU�zl�C�S�B����l��~E�]&bDR�N@�.Կ��XR�hxN�?H��B}}-���E��,	�[�3��p$u����3hBp����f`?�0�Tm�������10���Rxh{Ir|=(�x�#_�*O��E�j��ώ�/���rx��XĊ<@�O��Q��Y4R4#�p���BxT	�cLĒ�-*�j��,T�������:K���>	D�$��^G"���z �D�jj���I�@�`�i�N8X*�E8I��'Q��^u��@���.,�.�i=�����w���A�_#�N�*��ٹŖ��J������o+��Go'�AVɖ��~�c�7�~M��49X+Z�ݜ��j�;�=}R#n�[���k���}���M����Җ�q6$)U[f�|Q�<��$`#W��.�fh"jKG��ĈE��'Td�F�NS�� V3�pEv0�Rn9S�8C��;��_�����	�XZ�48�3�Īn��-�l�Eq�uM���=���{�黆?��R��-]���hwc�n�����᜚Sφ���q�2R'W�}���	��D�9��f��M����2t�m�7Kc�.�3^id�k@d*��n�#��?�����/J�� ~�	�2�����-��6���(r�W���8�]a���^�W5�JP����t�=r�ڋ�"á8R���k���}am�b�m��<]��>��H�S7k�Y�G1ڃ����)mNW���[	���G�k�'p'`���5gT�
X���X�O��!���hN�&ӄr���j�h��U\I��������;�H�$��v��9�Md|A�{y���S�K_/�G�f^쨁����*!s�8#�l�x��
:㋃Z���E�GB�U��j�:l[�	���G�������ȺL�?��؉3�|%�"K�yqS�.�yF�AT�.�(�$.ڌOS��U"Lc'k�"H���ۇ��I��(�w ��_J���u��7r+��!��}J)ץ���?IW�J2-̵hM���ֺ�V7���#χm�<���P/�H��>6<+�4�S赧�n>TG4W��u-C\��X��d�#����4` �(:)Lk"��P������P�J����.u��b�7�{�7���l�@�+C��%	
��4c�KZ^��8��i%��n��mM���w��R0=��`(X�FE(x���|�s�+U�e�>��U�r�{�j�鍄�����]�J�K�G\�U���ZM�Ym�Yt���&U�QL�5w:�<)�����0�&�Dz�¸���i�P�Z�v?w����:v&��;�zkP
���)�Ԡ�w;�`��	��+"$�����\�Y�&����u鎷ˬ��>�վ��hFƯy���&\JlI��Iw�qu�f%�5���O-i�z3��1�J2��;��%�5gl!޴�Ÿ�<�֎�gP�ZÓՐQ�}��D�b�|bR8�Yt��n�̅.+* �XW�@�cR�P��%�G<=�_$\�^z�ZZ�)چ���0j?�AoO����S�f<V����^U���v�Z�簟#}!����<��BU��k�s֚;����ǫGos�h�f��w����-Ȃy|��7��n՚��g�F�9K\����۟�m� EN��ꄹ�#��b>vx�����#��,��/=��St��lWUW8���0w�S�@(��.�L	��̃F7W�7�\/j����R2��|����M ��lU��/�Qd"Ga�Ѫ�+�c6[��^龿��.@Ai4'{�1�bHQ|�[��.zYH���Q�Id::��4~8͋��L{.1����r�*�",V(P�S��ҘKu"��]��Rg������bm�0㍦��<�h��z,F�|@�H'ƙ�KE-��m���92M�V!L�+�9�n����IM�N	2�c�1yj�>���(y����I�0�W���RO���.����^<�e�F� u�ȔM�MJ�{�޼�9�#�4�s�g�c9Pa��r��:cY�]����ٹj��"�"d�t� ��눛��Km��~��t�ꗬM�JD�l�ʂh�/����KvV�c���-_7�ω���;e��d���4��D/)[��
�B �%4�;g��Q�y����8m0Ec=�r9��/�9�۾�8�tXP~��i�h^�"��2�0��j��i�4�&o����8�+0�(k`�g��K-���bs�H8x6 EO�A��ԍ����c("��F��~$oy}z1e�v���� \]���]9z��z1��<s�m���4�h�~CmXs�Fgܾ\��v���C�ӠI?��3�W�ou���^H���.���0[�������I�&9����Q4��ʉ���W@�eB������GMf�I�t�~}s���A�W�aY�.�������zWO��-h�(s��wK������I8S �����q�Ϗ+A����ws������[�#�ۃ������;�&�V�*-�i�j� .ΝgJF=s��trɸ�ΌI�='�������
�4o�,4� ��z3�l9�	/��N�Hr�=�J�],���@��"��t3J�_��et��0j���4c��ɦ��e ���7d����V�f�缄�f��9
R������Gp��E�u���z�
��oN��TC6 �j`�I��d���ڌ��@���
���V�"8��/ �P_�RK�"-9�?��Gh��v���[8`l/�q*ح�jV�w��Y�i ���f`��c��B_S��;=0� Pp��$���ڜ��V��9�B#�g��
:M�{ <v�5G�靪�X�ٯ�����fQ��[����LϐE@̿z��(��1̨ެ�2�ԟ���%�E�{?��}���q��F�* ��U��9?X�7�����e1������a�������|�J��:���z44���U?�N�R�0%�KGޥ;�Q$�aӮ����B��w�fMz��,]]to�'\�����kb�����Or��.��r�����4H��;�R�^L���f�.�h׷��ȴ�
Rq�O�{���h,Y��Zm�Ϯ�[�x�e�н���h�wn~�J���ϫ��m�i��<���+f۩�����q���%[$��*��%4�18}\�>`�cp�֣yWb��l�1u�/`͐����w�ǆ����)��)Q��
Q<o�:M2QR��졸�3�k]zK��]��i("��Y��L4��+D"��o`yЦ��TLs�wx�ٖ��<n9��v�C�}6��n\{�%޳Q^?^�!B���.Tf�x6�h�C��J��	�hD����>����]��躱h��Dt:�qD~[��g��BR�;1����a��&Iouʪ��G��o���� ��Tss�4���8z6Ό��f�)y��i��뵴���WB>H�_@J�9:�-���MCN�@h)r���i��l��p�aܰ����O]i�~HBW�M��X��dM{w߃]��oك3�:�f�����O�B�KZ>����m�}�8R��	��v�<�M�]���� {�'�Y��@�<��T#�!��Q���?���q��C�U�I��)*� p�\+����^a����۵+2�eX ��U��Kr��E��Ę$�;U����BrA�ɥ*%D��a�c�oNx�I���:�\
�%�ܢj�h�m���I�mE��D�$@��'Ziݢd�~�!�A�@�&��f� �VS�a��Ā}��z��S�_BnU�������V%I;Z�v�����iyTǘQ�3}�#[yLv��@K9���\��J#��W.dv�s��Ѣ��+L�z��!�`�Bu�!���(��iV��;����F���|����Y��\�3a������Y�d� f���s:�|ߤRH�%�,@��^�.�j������Cn ��#,Tm:ـo`���}�T,����37O��JE����/� =�EXѣ�6{\L�]B�����p�|p�΋ ـռ��~*M����i[J�������}�_ �g���ۈ�xh���*g��w����9N��pةG�E0j��g�>Māu�/~A�d�)��"���zz2��#�^�R����9G�%��c�V�iR����S���g�7�f�z�J��6��x�.cb,�?�Ec��8,��o1+��w��͂��Q���w@��֭����a���
+���R��k:�ITӊ_�%J��k%N!NV�����&��l���l,`���u+�	�{>K!oێ{4�F��S^�����Amw"�%�1��bB�	K��Wlpڬy�@�1c=���*ֲpO�s ?�{n���b,����c�+�_��@�]0��95�.Z=�Ict�e�f�P1��Wr��`�(��}
�o��S����"���YLX��F �^̤�P��'�����c�E���p�*�GbYo!A����$fO�us8�c�cw������E:~x�$��M
���(	��ϴ�~�����-�,�(E�3�T�+�n��+����� �T��.�3GB���&�`]�V�u�_RT��|��K5��(%#��v��Kz�����Hg8���o���g��`ᔭm��Gkš�x�!u=v�!�ǻQ��#O�M_����U	۪t)y��y��
�� 9,iV�$h��W�QrI��#Ģ��|���	�ne#��-V*���8(�����P����a���
y_���{{/fR^�nk�<�!� ���\��wN	Q8k?�t1��z���h�lH�$���f���xO�.�0�bjy'w�q`�|G<�ڍb�%��n]d2��{�rk��O�$��oX��f� Y1�S䁅�G���Qrٝ����U9h+K��-g
��%��US��Fc8���;�%���\��O2 �{l���|��Xt{*�D�o
8�?6Q��v��;pPR��������0u뉔�ڪ�Z�ɀ2m�gK�_0�楔z�jϟ���q�ׇ��Ye;-CR��晻��%<��
h~� .�ޅȶ~l�1	ͥ�!=d�#�E�1�+7S�xwf^�m�2�w��2����8gtU\��^��+C��o��I�][nݪ;�)d�	�K�%s�_��%����]���ݑ�ײ#^N��r�_�h��C��Y�'#��?�Pj��t��8H�ioU{����N��Ǽ=��%��*��j@�y�I�Ȋ��_�I�է�я�eK�;�y���0-��+��q=�\��
jsNp�
.8���¬֒.�ra͓$��e)e��� >:��LБ���-M���s�V'��:���-W�l7���e��sIH�t�J�>�֓�y�3	�{l��P�SOt�[�]˿es���[7`��(@-�QEԸT��@K`&�O%=����Y�DF��� "��:����L�5���j����'�����ф��=�11�����=:3 ��_�K?���D���\c�Vy&��_�}ͶC�.$yq�;eՙ/���m��Ns��%��wILF,p�2�����;ql����G��zJ�l�e�{�{���+~ʞ�]��j���]�sk��n#N)4`�GlB`��ԨW�,JeWe�輵��^�
U����m�5S�k�d�NCEvQ��(�ҩkd�[[ԋ��WJ>�g��3F�xǣ3�{!���o�W-`�*�c���B=6�8�\�L�����&@p��x���Y��D�9��!!p�\�T�"�r����!kZ�|T�Rm��BB8A��*'>��ٸ�U��DPd�7<'D����c���%���J?�$"`����,��� ZK�ʭ���)�@���v{?�Ud	�P,c硑�������>��<MͰ����@zj�}�]J����<*�%��;8���������i��y`b�I�-�ɭ��{i�DF\ em��ѳ�P�ݜ/�(԰��JP1Z7sɻ�i����(y�y�Of�Ea��.g[��Q�����6��<�+�2��^��z���uMBӒc4P^n��Z��ۛ.eD1�9��W3Y��}�6���C����a�/������p>��%�S�/jd�1�'K�JJh~�0sv�j�3�ILLL���囻eN�vz��l� ,�7|^�z�Qς��$�8����ݾܨUf�8u���=���ľ��'F[�����%��\%�w���[�/���7��!k����h˒��֭��b���	:���b�|�<|s�q��
����}�[W"�ԩ��*-X˛�{����¸dQ��� N����W����>c5;�d�M�E�W᳛�k��|���'�h�Ȩ�*�/{/��>|j��k�0,�
�jy�d�I�`�N6w�a����h�]�XO ����cx�X������՜���R_���j3�K�2�X���,�3*�9�9��{�[Kϻ� 3�c�����0�N辬i�d��-fL��)ņ̘��rR�u޽�'+�6�Z�j93TwM�ŴHP)���(�%fp�ݦ�F��^h��#u���b�� �	��!�SӞ_>�<׊������W9��u��_�����ح'�5��n��ﰐQ�e�6i�0�j��u����T�������B�����{ݟ�e*�sY�= ĥ�˝�,[(=X��5ʓC�&@�]�B�;�g4���� �]�5������O�B� �x�]�����@��;ĳ��Z|��I1�ך�d�+���0SZ��o�{�u��)Ø��gT���I<��)���T��GҀJ	��d�_�!;��vn�>� �V���(+�s"�3u���m<K����f�~8��h��Ā�m��d���&Ne��
���U��Y.��IH(|A��I��#�m[Ps�TYA������+6eI�ǃ��<4�����"(�G'�D�ɩ2�9����,����Y]��e����L�ds�G��4��e"R�5X�56�E����}�ax,���,�О0�%�X	��I���+�4��O��� =s!�J�P7y/�	ߖ�(e����'T_���.t�V	��Ƞ�w��|aNZ�n6�kCQ7���� �q�(_�)�7����|$���A��M��k3��Fٌi5;�I����K�2�Z�w�E����*����t7���s8Z�D�RI̬�L�8�����L�-�1��Su���X>�G����AA��ѯ>2���n�)�^�E0|�fR0�1NЂ�茣��.�nd/�:��{�bKte�f����x�H�YBq8�F�4�������N�Tv�ʰ�ѳ;.�eZu��ff0_��?$H\%�����6��
�&>��%�����@?��r����x��n�U��}�C���3��ѽf�Kv�����lV�}�}+m)�|��I�9ac4y�R>u[u���aY_�����].e���DsV &y�X�Z��51]x߭"ϒϼ ��ec���P�U�%-�7JY��]�>h̉�M	���[?{�r�#h\�>�2�.Q�N�ݢ�U�J??�>m�!n�B�,��e�(�&�S��d^(���OoQ�P�����~�0�QE�K��Ny�96출�ߨ��R���n��K	1��g^��D3��G�k_��`N�ʗ���2m�A$T�}��|ljR�?�N��������C��}�I� ��l�|.D�Z>۸�Oɲش�s@���i���ր{��1Ӛ��8ɰ�� ;C@��a5L.W�^D���/���>Ѧy��HH[���bz��%�%k�gx�=�M���u�#���I����D>�+}ic��t�E����d%��_δ[٠ւ~Β�FF��6�����ψ9�9M���ŏ3�/�F-*Y�^TSn�NN���5C]�ٴE�$��vOI�uY�-a�"G��?��O����(�<�&�B�[nO��%h�G�����ܦ^��/�/��:�����j�դFʟ�cl�c:E�S�_-��ɻ�h����d[���)���y�#I��)N��Ǖ�����]�ק��+R[�4r�] ���F����jӓ�!��|����J�N%�������Z����o<*�
�ҿ�{! �O�	so�Jr�mN��Qrj� �
��Ғu3������~�'�
������N��$JCrw�1��$Q[�չ�n��2&�NGg??����(I����A�gWP�mH�B�!@d��+��#�T�"�gu$�N|��^��mD �LQ��)�v"�}��ofѶ۰�2hw������	;�=����f�=���H���B��a�*-WQ�[�c��]�3�|+t2�q�1%T�P�U�⅄'q�E��!��PΖdё��a��^Xk;�>G�sFH�e��lJ�	s���}>tƲ�����g�(=x��V6B2@Y
#�R�@-	?�d�U(��X�PV��Y"o96�6��4dϔ۳"�0xz�|q.�a����t����&d�k�+J��6�@���`v�pm+�o����%o�it�Vw>
ZS
5�Q�]r�Ӄ�Ci5�������{�w3�'�l���q�̏94��6���i�ק
�+1掠�L�L�=K|4E�dǂ���dËsF� i��_d
��%w��"���Py_#�VZm�\�y�Q-�F�����M�� ��9�!�T$�IW���>�:^��QR��W�^~� E~�n�EPt>��m�Q�u���/?h;��	C�HF�'�݂�Բ0Syjq��G�ܲ��`�:��j��H��X�I���:����;�����W��jDi�c/�����eG �?��� �����e��,����
��U��c��f�x��h�HZ�ܲRw�$����A�/z�H��c�X���_�
Lse��"��y>\{/�I<���WoC��9��%�,mz�r���(�$�9(�$H�ì.e�f=|z���M�EE���m�G_��ji�	DDQ���7��
Ϲ`��/�"��y.������Xv�s-�r��G�2��1��r0a%��2ZY���:�I�CuK8�hs����yb�ϛײ�'���5!m!=_�d5���� ���lX�+��]\�R��`���P����'0ٝ7�ޭ�GQ&�}�.G^��vch�p��y�B@�Waѡ�>�!aE���,���hP�b4���l�I�Sg�Ι��߹AC�񍇷�g��m���/6>7��Eҿ��}�ce�!�:<&
��_?C��<�S��΢"*������v�;ŋ���H:��nX�o8`4���uX�,���V)U�&2N��x�Qa
Q�.�Uf����:?�L�o���~�V���/��\������-i�� ^�R��4�fܝ�R��,���J�����x��U��L�<���9�.�;f���G=8�%c���:�u�����8/f�VK�{R�~�hc6��PY������r�K�7�ES]1/��:�y�0	'b��2���;SJ�R�9������	P8M'Bݩ�.G�4���b~���o�I]�``	���=�^���fq�A�L~�l��x���Ĳ��,�U�d?�(�@A�!�|y&f�tE�w�w��` �����O�C�ʽT:�� W����&�t����6����3��u�?tΠ�˪�ZV����^q�Ȼ/��?r9}�]+�Y���S��#vq�E[I=�;rc�R��JTf'z]����q�� .��s���Z�#��<)���F���]���K���
 8����ۇ�r�����2��F����$�!Kb]�����LgE�j�L�{�xh�c�T;1������V��aؼ{����g�J�%]Y���ksR��p$[��_Z�	�ظMˎ_��3��AԊ�}�R�h�l�z����0نQ���Ԁ�p6��/�z�VaLBe����.�v�RX��F�G�^K���{*HR��⳯��V����cX��QV4l�1�Z�&��:.f��3��y��ܩ��o����^9d��0�ޱ8V�����w:�$�͕]��� z�3hC��X� �|3Ȝ�cO��pf.�Ҥs��;U�5�@�#���QІ��H|�!��M�=?ӣ�&�` �Ij�@�Ѽz�B-��71��f�&9�n�$�����m�KT�9���'����qa�4�Iv��ā�2ѽ�z����*�~k����(�S�w�,݀\�x��ZA=5�պ�%DU�� j����4���'�ₜS{T��":�Ϡ�ȵгN$��nG�/F���#������O�Z��I��<��{���
q�!�Q��"��7b�?@�4dŅւ��=�)���y��~��9x�_ӥ,�:VU����$��K*���.Ң:��g\\HT�v��?���v5�(���+
-�����k���˝]��y�c�f�_�u����ͯ�a'�AW/f'D��Z7,$���^�Oؑ���(&�*c���~�ڮB���N��i�7�R8��������o�_z�kywa�t5�'�30aA�G'B���;vF?��U}k�籸�1��S���TJBk^�ă�ϼ���� ������9�;��̛��-M��y�Nu=iO�P6�nT��I�%�Y�\�+v��s�#V�����|o�ԫ�m*`�Z�F�o� B4
)�T��:\yH����~��,"�5���Z�S����L�,+��@x��`|����c��:u�I7f<��0V�,��=0bk�a��sl������ȓB����/�ǹ�N������Z�f+�:�f{>>�O�|���!���ў3��J�����Y�9��H0�N5����_���9N�K��<�55jX�<��J`��� h�ێlC��n	�s6�������0N	]uV�*�M�����v�0L�I�7���o1s�S����2w�rt��IQVċfXȋ�L1�L��z�[��O�0�Ω�s���IT�[ v�e�"��M�NR��p��B�:O�Ep/�kʾ�c^�U�~g���r�P��	�*J!�7Nw2����@k~���X6�=O@�VI�7-R�.n�� �Ob�������.-�)���� e��!Y�D�4�dw'�$m�L�zob�l�3���_7?xb�-°�zp�È����|#r&y��7)�����rJ{��۹u�ʗ��Q���lz^Y�I����{�{�C"�{θZ�Gڭ}��ԾT�̯R�4-cj�7ć�U}�rJE��[xd�m��]�U��&����N��9n��p��^՟B�c�=d)Q�w9�8y���9E'�1��O%���������Y�GH�ũ�w]YX ��"�Օh�l��-ꫠr���e�P}�#�p̕��5�uQ���Z-�r�h�SE��}_)���Û��:WR���}��3Hg��0�/)TL��Tg�P�����m��!���RP0�>z�Ռӎ�M�o
���;7�<��l*;�N'�"�e�G.�>�šݜ%����y-W����bg8 S�[��φ{�
`�^kO��a�#�eVX6�&�*����J�(-/�7f���γ�����UID�XҼN��!ޕ<�����]ұDe�;�\f��\ ��whd�<�&��K��x��	���M����H�\�w��� ��f)���+�����`��x�i���W�Hy����pI@.gŠ˅�,��ԃ�O^�=1�#7��2����_��7O7񔱆�]�P�T�PK��4a<i�&yo��OF�����1)��.�3����bz�:Ɉ�/R;�Md�J�$ub��`-9>��h��Z�%4�8������kuL3�Ȑ��xX�=ul�:%���t�%|0��6O6�}�A����ٳsh�.)0p��ˤ�V� ��i������Tw���,A�Xa�6�sRZ���K�K���	��R���G�_��.�t���=�6�nKC��i�u0�K��[BC1k:U����7e��|�^8����$B����\4��,���o	D́a��dD�v� ��O���I� ���@��C�K!sK�dK�vm��>5=�y�o���ߜ�iG<�U#mzߨ/ܻ�	��4J�3��:ͨ1?8���so_0��$����TǠx����:���E�����2����̃�98o����x�1
���p�m�Tnq~iU���8Q����T�����QDm���r�q���Hw߅:]5�ѭ���P�d#G��Eo;=�
�9��~R��]@��g�w£�Q4R6P7h#7i�n���t>f܋ �qLB���)����
*�U!���3���뉣�կ�
�6������9�7���#�JIeS&U�d��i�JB=\t��p��A�M	�'7��1��xV���H݀��U�{����"�=�/9�a��foty���Ð��ac��J�HB���X�Ȫ����:�)�|�Ta��g�m+�Ôճ�ɯH�v|��YL�[ލѨ�81� ����q�p<r�fvu�c3�����)P�Z����g��Q�&���Ay3�a�?��y-���<btzSb�p��sR�C����S�֏�02ْ����?�F�%;xѺ��hm3�˸X(�ΖU�#)�`XR����tCg�`eۉ�'h��r5!j�Ѫl�֎���gjE�1�';����A�R��@\c�^K"ϟ��b��,L(x)7:X������\����5��&|R��;���y����k�>v�����P���֟xɜ���r���De��4���v���<�?��~$�.��f�aؽ����Y��q1&�Deߡ/ g�Esy�~���@O��+��~��Pg�^�IY��L*�~���F[m���'�!�7��C�e��7���(�+P����O;��)��6)҃�_��Y��KP�%�1h�@i�2�#�ĳ�;2M8�3�
蓅����o�4��Ő���K[N�Z ��L����̕af��q�A��U�����,�(ƣ���
�,=��hd0����M l4;�a:cz��M^���s��<��~Z�j�DB

�}b�l1:�۝;�Y�a8=��VQ�Q���2 ���$������S�p�z�(y2"�>�W�)f�B��x("��
I��b�{�d7�\�3|yn��vd]{�Qi�j�iU{Y��sS29tH@�̐���lAIȭ�!�
��U&��;����E�|F�O��@؜����4��r�R뛂��@[���k$�W!:Ey�%�!�~�����O�
��2yu�#u`�si}ұ�R<E�o���E
�ctg���lL
���!_{�W?1<���C���]�~�uD�ytR�fm��2�!��g�GD�vN��䮜c"M����_����p�d'����������x�W�U#��P^�+��Ax�z�}ʄ�k�q�0M!f�7�KQ��Cy�U�8<u ���z�����:we�%C_�����zط��^��n������c]�tҢ
�,c�j����$���K�<H�P��l�u&i�(�zS�ГN
!�����D���!����ƫ9�bliX�rS�A�J套8X������p����o��n�o�,@�(�tܗHSpf�#��� 2Mq$g"C�R�!��<�o�X��F0MU�>�.�k]� _�w{�r�/w�y�W���,d ���E�4a��E;5��	�߆�@$�h��dt���8�LQ�8�D���4�Gu�'k�WJxF�n��=�.8������M�ӊO��m����䈺H�n�,z`뢷��G�V;�4�c�r�%t�G��b�����DK����3��g˰*���M�����m�l߳���Z���+����!��U��F����ʓL����Y;PЭLj�B��C@��A�����X�[�@y�T�D�KN�Lw�"<i8����B��?7_q��mB��m��:!߻��M/�&Fd�YfF8_����D%�;*7�4
�#|l�ܓ8��v�� ��F��f���V���5��a�f�����\� �A�z����?0�b^��͉�t��!�
L5!tJ�)b�l��7���x�����ɻ�`J����?�S�l� ��%Tٻ|�؟>��~���R'C����,]��cJ�m>���
P�h�=�_k�K�>�6mFu �_�;A��9I��+!��߃��Fqˈ�U/yjԕy?���eB�0�[���f���o�儼����90�Y,���57|��=;şp�I�����Z�L���lm�<3��#PE}����4@���4�05�BQ0E�M�`�g6��t�Y���'u�~l[���nZ[�&��i<���Z��m���$�-��FEe�	6����M���u>���?�A�p{(��2�k�rI}R2��A�Q���}�M�mL�j�SJʼ$ve�e�L�����j���6���o��U���+�;�����G�#(�*�Q�Q�QY8�����ZaTBT����k�v��dH
�*�/��/��2��X���X�B5�����G��];�W��l���At����9{��*���}+Ya@�&Z�o��+��.��G�y�`��7��dW;�$�����9����z!�sOY�yѼ	�o���%��^��"�/�����:��I���:��|��]���j!���q�ʽ�K�� )�]��F��g!Z,�6�D#1���i���������z)5�}{�U�_k�j:e��k�"juy�h��ݸ��8�K�:�kFF+���~:6��`I�ӡ���|6�E5�����i3��%�r�������OtA̅Η��H57g�w܌�¿~���R{���i3�u).g��3:�fT��3��ޛ.�Z��3PqƋ���p9m�>�X-�V�n�̼��y��0�C	�1� �F�mJL\`?e0#��5c����-�0L���`,W{�2�3�LKePM�����nZ�%&@���|��RE�=s��!�דq^�p�d�_q�)T���Ft�'(	�F��[T�G��)�j�d5�
]?�&f����Ҹ��.����m�q�-�����;X���@��B����:�#!T�E�d�����z���@�]���Lye��Вh��~�^����@l{oʷ0���hS�Dnf;�/�d緧N�ossm�}R���l�����D���$[[ �,J�[he�:z%���܋Q�?��}�&�sM�����MU�G�"���~sA6)�>�N�ʰb��U��Փ^����x(��:3�]�g�d�b�K܀:�\Y-'���w��'{:s�"�t�Qe�y�����&l��O4)��ΏLϓ�Q㛕P)_ܩ����`P�a2"'�Q~8�p�=v��L�˜�G��~�h׼��� �p�bdK��t�h�Q�g�3I��4㹮�P�.�t��O�˗t�_�$�ݥ�+i�m����F�LT@U����x��\Ė(B�w��J<	CK���w��˦ ��:`�Rj�:��߂\�^�A�[]�ٷ�b���ڜ8h�tc�[&�$1ݙ ,$�0<���e��XԄ����a|��H�vtb��y��h6/����,)^Ac�WE\w��Qv얶�_�EX�����m�MCH�.�ӜZzy�`ܐ/:-r<�1�0X�;��2N�0�D~�e�IS\�y��	���?��ޮ7�t{�c
k�q��φ#�Y�'T��Eja;�)`9�h�g��ޑiU:���=e�͗��� �
؜p�N�F���-��"$AL	_]�)�P`�KlM��ܒ��p����=Q%�Y@���%��'MmI���2I�)5��c��ɔ%<3F酚���з��a\ j�&<�r�$�<�owt��L�A���ps�ᝎ��d#g <$,0�v*��!��@aa�B��QD�ZM|��8�����U���YX�%�G��w�.����s�h�����n�ˈ�h
B<�r�����QV�E�s��l��l�k�Q�7O��w̻�>B�%p�ң��n=�@;�C��C�!��ST�d�2�*��j��n
��;��;�9x���:�Xڟ�8�n7;�r�v.����=>&Cw%�b	�X^�!NAw�*Z��&��0I2 uW+:4����c-��x�T:<����a�n*j�U�����L����A�
�<��q��Ld�R�Ӌ�P|�Q,�8丅9�`!����1��)Z0�U��N�UJ�f/�~jA�V����D��5��ERα�x�4E�m����ˉڃ8<�P�ꖒ�#��'λ�I���=�e�K��g�Jݵu�w�>����~��k��v�ʋ�!�)U�6p���cF�Єy�l拉��"�m+EȈ���B)�2g ��I.$���
v~��-����$7j4C�ЊB�1����;Uib�eC�����~��J�˩�ö+�.�#�螆��6�i
�&��|��)����(���9����h��P	5p�t�O���hSW��E_��U>�M!dO�:|�\�	�]��^*����"�U���׺��KZhaTx�G�{�U`���}+T�.�ڞ��g�f�f�oAIC��lJt�玻N'�ɂӯ������JK>����[�k�L
b�� ���-��{����P'�o�)0���z��FT��p��YN���T'-T�[�9�ۡ��Esf�L�i��O$�`A������
}&Z����tT�#��lzw��~� 7z]Ѥ�x𹫳��#=F3��d���1�\�L�gi���L�%��ň$�Lb��1�}<;ӛ�f�H=�
v���� >ֿE0ۦ�+��$1�M�A�����SQ��  �k#�Z��̳�9M&ӔR�ᷓE8�m�^f��z󺵠���~��.�����`�P��9}�J�����]?3��2E�RmV� f�5�1������M�������t -��N��-�,�0-�}\�����E�ۢuu1{�zU���H.��cJ�c���]�+>��؛�A�p~S��-5���֡�Zvr��4��+��O�U�~;��o���+�O5#�X�b�����E�2�4!�tu�<��$!���>>D�­B��|��;��f��`�d�0�TWc�)��>��tw���G,##.АJ���{��k������E��i.̍�S\j3�bƇY�76҂�Y%+ǿl���.��|:��jg��3����*��KGzi}����j!�O�=��T���d�uq*�{�t����>𺬅)�6�ܨ�\��\�k�Q���c'B���>�2��*I�O���A�Ma�V=�x,-&ũ:5ퟄ]~r��#��8e��?�"�����e[aB��伇��D�ϔi4�-5Q�0,����U'�
DLIu�n�&Zc/͞�E3�Uc�nܱ�pU�W��k	�̛�.��2ϛ-=P3ϴ�������jW�����j¸�͡ByRBG^K5��R�Y:7��	�wʞ��s8y�`�� �[�`�_$��S-ג�y<q\20���y����$��:/���p�;�eS���<%?p�=!��~��b��!��4G�+2�/\���"G�CL&e����ؓ��?��:gAd���7�0�^
�mz������/��6G!���/0[�]Z�É�G������øK����g����/Γ�d�!��\��B�\�W�.���ՠLWL����~- �[`��ڲ�U����O�\`�,�T��\`s�3mp�I�!j��"}w�R��.�=*N�G|N�Q�Cq]$pW����GbD�8�)_��^5A�n�"(|^hw�힣���eՕI�b��#��-�m�d��soe���n���P���JO��Lb��0N�Aތ;2�ԦuHI���9]��N̘��j&� �J�x*��խJv�A�S'˽aS�(7Ǧ��H}Wv�4�8�d�ϪL(�ID�&E�1�UkI��� ��e:�0��p�rH��|�Ʈ�?n'��1��wQB����$��r� �5���kų�f!�79M6;G�a'd�n�(��Z>�>&��� �w���7�9���zB�s���,٬���5RJ�3'����2���	Ag�Rߣ�6o��4�p!y [c�O����M�R#����̉��y�EF�ygP�5:��!��T'�J�KAh����&����ȫ������c�{�O�������}(r����������N�&@��y7�n'��VW��^K�u�	��!잠$2f��%u�+��M:vj{~`XZ�2b1 �t?�N#�!�.`���<��/5邒hv���z�q[�B.��Q���64z�m�*�������>B}~
#*�iC����Wv�ȟ/��Y��Q`���hJϙ���)~�gr�:�F)�<ߞ�'�G�4\�a܍��CDCƹ�B[����v��9Rt�w55�����I�QO�n�39r��\m'ʴo�6�6����w����ɳUͼ_�&[x��"a��I��ܴ5]HH�.!L츀�Z��i� �=��>�֤	G��ZA4 ���ڣ��H��+���7׶f�ͣ���g�g�+4��	�eL���-N�_�l���X|ӓ#�v+����x .��y�.~�ܞO�L�f̧ �D���N �P �R���O5��O,�Z�ܹp�0�����X\��Q�C��k�k/8(tS�]4���2��E���$}���l�P���'y1�����N�/a A�7�J�S�k�����੶��9��f'�����PJ.�a� �M3ĕ\����`�A�\1��j����l<���-g]��W�.#^�~ʁ�!�]'�W@�$1��%�2@�{��V�0R�U���a��͵h[bԖ�o�4ߦI@z�:�p����s*J�G�j�=�����آrz&#=����K���*#����IF��q���šd���h�Qm��Ŷ��>M���o.z�>��6��-FE�LkO���"�,��ｍ��0l[�m��*�k�����3�kA�ǘ.g��R�N���\��z?~"��3G�&�D����|"J�\��`�^���kCFz8���AcN�坄�$��0��>�7�bӋ�}�{�Ⱦ�c��T�6�4���'|Gx<$���)�P�+�����`bԒ�m�ΰ�'* �k:d�`P����"{�)m,�2�>9� &d%.�KoB4�  כ�� 0�4"7&i���=`~��J�ЕС3n��fw��{H0��P�xK���Q��&	�|�-x&b�;>xY2�0=����_	�i���g0��y������&<��/ג��=�n����<�7b lQT�C��q,tjf���FaY���GA׎��ey�pʂ�$eJ8~/��S0A����C�į�ocD	�P�\J���5%M`��_�kw7��:ɪF��\q�=��;���QRr��t��T��$��|Ĕ��,QՍ;"�����_WgΔh7��G	nQ	�ƓR��_-�E���o�e��7P�����']�^���B�>M9��z�_P�ET@X|,�e��%,�=Cj?����+W��F!��)֋i�5o�9:�}�.���W���bT�5x��ꬒ���B9���BLJ�4�=��˭����@���Gy�U0������O*ɩ3Dw����Ou���K�T\>pW���!��Q��ߠA��q�Q�S/bIPT��r�ׅԣ����ϸ� :��Ky��2J^��RtCLʇN�_���)Z�Fn7�T{�͗���^<
R�aʉ�*�w�n��֟r�1��T��L�y9��m�C����S���f#5�
��f�y[��SO��O����UE��@��.� _�y狣��v��$Ǡك�N�|2Bím�����s�i(�z�ˡ�Μ���F�*���������)�Z�8�6�=/0�;�f�~B�л-�g��{І� �z�X�^�u�-�OH�hʹjNB5:��S`��[���'hi�	� \�����Ց���J��r�t ��q�P�TT%q>�n��h�:������g�嘞�-����>�Fc�k���ʆ'^Dc�Dŀ=S�7j$VF·�	7�sC��nT.�	z

�[v��� ��d��'2�K0��>�k��Ɓ�Ü'��ϲ��N��f���}ڈ������,��d�9��q��1�pl�ڟvzk�<
�M�����ZW��J�,�8��(mt
�@�El�"~�K�`�|��ʒ��>am1Z7~h�o����2 ��F���H)�t�٧�n�N��]R��� s����l�#��� �M5Yg
��c�&~����2�Sn����;�֤�E�_%)8�J$_��Wyg����wDo�ʖ_���y�KG�1	�E�qrI�_�h���X)8=��K��#���B�q����#k�V6W����rIհG�G�j�7����II�xT��Y��)��M�����i*�yP�wQ(�ۅ�vi�%v}iJB�v��;���G�mG�P�?'����(߿R1�,�ҍ�X���[}��A�O8�������DQQ�h��U�jM���J	���"�x�M�`�,�Yr˛՘�[��m�8廷��D�̀�"v�f�[��ӣ�p�㫪�9.��=v6�/�1/����v��]J虄2�%�ǐ�r k��ܼ���o���ȓd�	6d�U��{�rhs�`t�4��h�Yb(w�uϫ�5�ȭ��%3_62��1���R���X:o#Y.I��35B;>&*�Ӫul��b���ٮ�f��MCI}���\/����W�d[\/��Ԓ�Ib���r`.�����S�l";����TS��.�֡^�5�a!������4n�ݙ��l��ffR���xM:!���	_D�8�B�e?:RB��}Hh� o�q�42P���N�׬Q՚�j�U6]_�p9�/����b���t������ǡM����$R��!��5�~{I	��s"6ad���gXj�)^+�Hcx����{�g���o��t[�<�
ײЯ�������i�����Ð�h���?��ٌ!�ܹiu��q��(��Ɖ�q(�9񃛄����w�s�6����ԉ1uU^�K��p�	�n?7<��`o�18�,�y�Ё�����p�_@
b#ݕ��������!�f��>N:��\;����}�#�M���Eн�Ӊ��t�x��h",̐�7�E�p�ҝU�%�r�WB�}V|g��4K0%A�И�}�H�����F���t���a�E����:�mJU@������D&&��˫Y#�c���ʛ�w�Vᾤ�=Ou��U�ۤ�K3no*֮S�g ß~7�,��T;�p�6��h���VZ�DE#�ham�r�H��tA&SX�
7\k���4�O��2�� �E
��	�q��R���\~��n3���t	�u��Wn�%�z� �4���zA�c8����&����|��r��I�x��<��T�W��p��Fd8.�2�Җ��L�tq�6Z�ʙ���Y�#|��Z.#��տ�C��YB����Ke���W{��;��I��<;c�Bjz�<��O������t�C����$7n.�y�D�����s�� �J���q��Eo~qR�W$ފC�F��=��42a~�`T��g�hfN� ��M{��.�3+��!����S�>��o�J��p��yJ��S�RBx�ղ�u*6PR�垩<��Rn�a��>=i�0�ۙ�PMgC����V��V f�橼��W�KA�����*J�[�Jel��k%}��%����vU�=�a����C�LE���V�.�����B�FF������n-�k�����Y� 3t���0��\�`�&��>����BibI�!ݖ<!n�OCUJ��W�Q�K�Y���LoP�,X�4I�zW�wx�� h�n$q�P�f(�t(�2�5�����{K;UJ�t��n�E���h�$+ϫ�47�`�:����l�'�▿�i�.ȓ��� }n�|�*�^�h��~Ƭ�-+�`!�]M��@G�� ����1t������<���4o�}�!�z����8�cY?�|�]����6_����a(�t[!B�s��sK��9�l���o16y�Z������Z'mgLp���T �ݛ�B�r�@�qtO��o��b�͏f"���ۖ�N$�dˊrE'T�<n����s3��Um ���cQ�=x��be��=���G��m�!\"�=-�����|oS�At8�젉0v*S(�9�>UT+�B�Ka�d�M�);�E��S?���[g
�|��i��_���ۇ�J
Oa%W(Ý�B�f���?kB�/jq�M��9��^wF���JE�����sF��H��Ճz�qqbM�0E��d���ʪM���I�}�����G3�"R�X�OJ7��ҺoM�����״�\~�K��
k;B�V���2�r�JC�gȯ�Գ��~84�(��n��B_5,\f.x�����o ��TQ�?wƶ�K���DguN=;ۀ�Г�q�����o���3K]W�/�e������
�M��h�/����󛟐T� ݃Wg;邿?�Ǐ_��)a�����}x��W��L����
��S�gyc���$����S�z�j~�f��c@�X����j[ �Ie?��Z�� �#�w	��^ɨ3&��(uv�-)�)q_���|�� ȿ��b}�"lؼ�c����JJ�͊���e� ����Di�F�oș�o�3c��%�`8¼����*��|�\�������-��=�D�Hry@��3�wB���WJ�l�qi�����j���F��%Lخ�Xر^N��ĭ��c?��+�a��[<��|���۰Dv�� y��@���QD��X�w]G����~%0͔K��� ?щ�lP��yC:�q�g�V��w�k�x��������ǫd��O`åA␏�bj�~��Xb0��h�x�C�F�)�y��|}>���Y�?,d��d�����3{�:�*��i/�`��m����6��B�ڰa���[O㽧d�|0�C�$��M)@uDo�z�wʺ;
�©�ZL���P�
��d�D�³f��d��Q��v]�7�E�GJ��WFd�R�#$5����
��$���d��*e����'�j`�d0��X��B��L=���aM��Ҫ8�*!S�S	�ۏ�3H�x�D��|�S��(��+��
�"/��=Y�^�^��LWNkg^Bd0�5�\�6����l_�v;��phL��)�2�璈_�w�y �nd?dU��s���	,7]0�h�*I�R��_��� r���>���ʎ��s$�[n�4]���^8���A��G�u��Ćԇ��E�n��&JZ>Q��13��8k��ˮ�	#`����U��'1�b�q4ۤGDma�#��ٮ�$��3����_&�Ztצ�c�B=(�[��ވ��I ��_����*Q+�<��G%_��ӷ��G�QC|f�j������qGfJ�+9�1����W�6�3����'���V�AC�ۦ��$4��z�z���!ȳ��
�Z.���>��U�ݷ���0t'��]���	�A�r��f�#d�K�Fs�l3���bT6����2���=�wc��$�'�\8@#���93lŒ>D7@�dϻh:����Q|~#e�H�`�f��W^���!��F'HKD��v����a�����(a���̝�y�;��(-��0�!�{�/��φ�lP��U#&�'�7�B�Eáh45tP��ɹ��Wl�Kv���3��h+�"���
BN�p�GKR��O�>,�A
u6����8da�E��ю �c�*�������T�,�����Ȕ	�����n�0�J��'o��-�������۱�@�Y�Y�x����NE��7(������.w�$��7�-��s���	�c0�-[!?� ��-���=M. ����h,feP<����	�;���I�tB:õq���u���4b�9��n�I�V(́�j���N���`ֱG�لz�ʁ5�i���z�<E��:2���j�\4DY�sأ���>w��Xՙ��XٱVG\�ҙ��xz�)��^Y\����UUf4��bl��Fc�f���/­��쩏�]3^���Y��7�6+W��s�,R>���SB< �Xƀ�iH��1���o)h0�N �+&>
k����@����$�gЫ��%Q�ޱ5�*�P����<�X����e}�tw�,}���r�Gf�N͵LR)��
DǮ45U|�`d��(�O-qu�}/�\?W+���rz��S��'5sL��˱@\ʷ�j�6Ye�S���'g1m=�
L��K^���XA�2�}'�/��d\|����.�肉(�x�6dnL��������(��X��� t��ɻ��f��iI�ʭ�M���`��T���_��вy�UOu"�۵�(#�T_�V|<r�D��lt;H*E+���^rcF�[�tF99�q�s�@�j��N�G�-�.�@?q�@ ������=���dŋ�a!�&��\A��M�\<�%�O?Z�d,����8�V��r�\��y�w�o���~d~��h1��&�"��~Ҫ�7���;� ��'AD�FR��V����Q���4,�M��F�"�J��N{:(�����=Vf~`���X+�^{����$���2	�E��Fی���[SE=QKH��E�} �1����xObkWk����V�a@�uV��MZ9��]�Z���w��-�~ �L}�N��!T�.>X�7�Gz��Xsv���"n��(
n���Zf�[L�Վ���9�|��5l�,z#���M S�4��p��}h��=���,'�gƿ��
;�@+�A�Ex(D�rFg���{�)O�`3��|�)*O��qcR{m�����H_t�*��_��>PE���I��� ��*��I�[�����73*"N2���,��]e6J�b��m���<�����=T˚~�>\�cY֙����"�o�J������:�����x�c������4)n�_M��CP�y�_�Gćȅ;�������{%�Q���C�1�a�����V~�=�Y(0J�֦�B�V3�ٳ3�X���o��8���pԉ�Y��JhzX�@?���\5�E�9�D�寶i�X�K	׮x�1���w�j��wͺ�b��b6K�÷�`Q��s��鄿�?K�{+�����z?�Z�I�*`J�RU}|�]�p�M)�A���7e<P���7�v��c� ��X;�����Hm��mt�5�b*�L�5{xt#��:AF�V���/�^{���@���3��IY��+�?5��=�a�C��X�鿊�U�,H��wt
c��5,��aRI&�Lk��y���_J��:������-�E1�G��T>����ְ�C���X����>h��=[$�*j����D�U�O��o��z�n�03AhNs�hw�D��"ԥ�1�h�GĴ*wm�3��_����`�q����f��w|�A��r�C���D@I�e�t�ny�(h*-̟��&���Ij�Ӽ�{E"�&Z�;�6.B�+%�V��2�����)�U�ꂧ�xX��8S�No*�s��KD2#�}�$ԃVB�ه��Tӓ�/�@͇�Ϙ�DC��o�,�-�V��Y�e�y�%���9%�=�9�[b�1	��!�ᷘ��a;���i*�̾ݞ�WN>c�����o�6�)1�~���$�|f�A:"��a�M<E�F���:�o�4�Y���`��>�|��`a7�0��RM!��<�¨𲚖����c`F�Z�I�O� ��t�2�䁺�e�s�Z�_L�U�ԯ��Z��/d����K"y�Q�2�Ic|�J�NOS5����/��E�C�}gzJP;����&� �-����C��M)�%�?X�1T�"ٱң�c���|c7-�7�2�d<�tBs��х���X-�u��DNk	v��cQ�/-(����Ki�u(>��~z�呢(�]b�Gظ���P�E	(L�|Q�j`�&z��0Ur���e�� �YՖ�Y̅)�2��}��+�̥��|���դ��OH���T�`�z��C�f��{�O��s7"b.�����<���ݪj=���3Z{9�Q�',oj5�o��_F�\U}���F���f��D1uWO�7����C�y���f�H:���3 ����{lYD��·��ໄ��rt�-j�� h�r�Vf2�\���R��H<�.�	�e>�Y��M�ls8��9Tؖ'ɓ��w-/�C@#�ނ�-0c�|������bÇ��l�����r)d*���^w}G}���ڟ�L/�^�!i�w�ak!�L�,ڱ��j�����:}��3�'�C]⺩5�s���9�E�|ݜ�F�6�G��?��Ǐ�sb�J<l@j<��b)؛�쎿��L@����_d�)��<nav�_M�sp����
1���r3fOj��~�\i�x9�,l�,ǝ'Ks3����b����������6\��Tn���{'1-����7آp��c�7iC� �8a�_	B<�V��Bs�"_��f�Ҽ+±:X�TFN�͵��y��Ak�J�@�U�����n���X�e�$֫H��o��W�r��a}QҚP����T��	��̋3v"����*Tj+ ��^xLu1+����E�:�>7n�=��z�.ߚma�q#�,����KU歝��I��>2��2��7�/P���C6\�����oV,h2�ȋ9��?��$#�r/zI�D_��5�|�xr�l;5�B�$��G�\�jM�{�j�b?jM���*bޱ�5�~cF�mvخ�����+����=Y��2�p9}�I���I�4Ѫ0w%߄��3��/�,�X^g�I���;3{���ƿx1�5i��-�N�)��:����:bB���h���u'�UE�P3`���c���Aǫ0��$��[w̑�4�*�/ׂ^�+�	3i3͒Hې�0�x���m��<C��'a:#�0eI��0��|��D:Q�T{Pؿ��vҴ3_?פT^�l �Ď.��R ҿ�̮l ��H��ۅ2*�Ic��`��+ͺ���Y��O��0)B�Dł��ɩ��;�8>]!|{n~&u�k/	(��kO3{=*Iؔub�?��R�(an����gT+2��.�R�TO:��e�9���|#�0��Z�m��U�q�(`�nW�C�3Լ����T6=}�|�6�'7�M⹿���Ke��}S�_ͻ^BsK�aY����)*����H�e��v��3��j<u�d�����5u�����+�,wW/�<�2b_"�?��O�Z�jm���E��N֫�[ڈ'?g$���_�ǖ�Cm��T��Y�h��1�����)�[h���1�rܹG�#���MA0םA��xK�W�W8h��9u���谘��t���X)�Z�MY���aS�~�3����%\��?MܢL�+�b��_p�f�1,'�������=��x�|��t���W��	�9�k�l�6Opfʌ�J;l��@��l57�����{�#y\1��'�۪���^�9��P7-n�X�;�DL�:�2٧i�V�o"wĀ�NU9�?��s ��N��VOk�Mt��(���B�퓒�³7��q���p:� ��TVT@2��q�33��A��kȠ�*�X�/ݞ	�E��z�ɻB�m�jT�
Ԙ���.�ٛJS.bEaZ� tc:(�&.�����m���|'�[��e�룹\��o� �Q^���1����M�'⦳#�x�L�j�S��gA��H�g��>d�z=ǳ�
<��x�Ҁ��t���N�tфh�^W�\��+(��C ;�Ų��Zu���B>E&���z�GyI
��n�O?ә��+[͎�&��.�2#MU�V�����.����Ϫ/��$%%�Q��(A:G@��Z�d��hӧ��9룮�6��m���6�����j	�]*���k�\����e�w�.���
�6�y����O/�ȱL�+�Q��G���7A�V��{��q���8��]�dy%ɠ�~Hvg'��� ���V'4^�~��{�w�,q��:/*�&�|���1�Һ˭}c5���~�M�F�q�+�!�t�K�E�T��>k�^�  ctFKDH t5���� �N��a����/-r쁃'D'�w�B[�Zv�6e/'MHIXg"K5=E	w�kʒk�F�`���`)��Q����
�4b�{ߤ����ۊBAC�z�!�*B��U��IP��F)�6�Z�E/�}�#E���Z�h�S��m���7���|SY�kC�	�����e�0��]����W��g�M�1�(H͚ذ��:9����d�!�����%Qv�i��?�b�"w��f���`=@��d�I�x���r+l�n���B��o�d�)0@���i�(/:o5ņG�97�e����3�El]����MO���n�,UD�;��04:��D�sUxޕ�F>��2�(�sӗn����R�{(�G.l@�4��d�C�]�7=�\�Ǒv���9��6D%�>Sz88q,��و��@@{���r�/oф�e����+����?����R"S�4�!�O���2B�c�qs�"\>��dV ��A,��h��8�?q��m'��8'2g{�&��Hj�'���zv	�3�F������"���2�΂�H����^���[�o�����?1�<���e��E����!�w��p�	p�{��Vdx?���6ȋ���h��@�+�E�m����;��F�Z��͙�=gaN"�Ph7d1 �fF��E����NNQ���s�F"ծ�v=v�1��%3#e�T}�-̘3�����zϱ{�=�����2.j�}a�O��]�I�Nl�DB6�w��_�W�v�����!P�tN.W�� N�k�<[����2%6i��z��i�h��S�sn���E���n�m���D���ب���>~�cm��T%����F��ኂ�v?}P�J���i�)yZ���M�+O�ze�0ຊ����Ȧ�Қ�X'�32ȸ�}!��/yør���ش�* �Dۀ�T����ܣ�f��7�_�M2�M{'����@��/�a�S$��*._Iu��� e����K��D1Ug?��/�aYD�f��Ay�ȧ{+p��y�������@�kt�t��~��J
�e�]�*�,<G��1�z�����Y��Z*U>��� v�p��Cz�H�e>�`�;��Pr�;nl��ȸ��p5����+�[̏tf1���pɇ��UQu�_�ۻ+iEM�7����W��71��?���^t�^�,t�FJ�;An�8	���3�|ow*LB,�M�Fr���S�fJ�%#lD/����8E����^��l��-RQ�BA1hD}n>�9�ٕ���yhcS~���Fϕ9��pJ�;�<�]NL�:������D�_PI�Ge0ó`-^�_�_��>&�~K�V]	���]�Z$��xf��f?���Wd��-&�{�l+6�O�%�j6�B㝸�d P��΂u�{�4"��M��ޓ�=�⇔6� �!̻̖Z=h����ЃRFir��i��v���&� ��0<��s���bѩ���a�h��ݐ-�r	��nA�%>!e��>%�!�����ґ!����ꅃ��W���qq�A��f|B�?w۫2�!��E����1[=A�M��Zl��k��ݶ��>m(���
?e����ܾ�Fr�G�D��x1L����h=}(�cet�>�����窎���W&Z��xH�_-5�`�yl%���2�|��b{sw+2of��Y�E����t�������3;�=���/��M��t����/���	�81'�FJ�cdڹ�ѳ��[Ğ1��0��Q?�-W��-o,c�o¯B��25g>2�~�jAГ�C�>�
�>�ë�YʞvP����z������*��Ɏ�O*!��v-����Q�j�)'�*!�˦��_�*��z��b�l@͎��4��?�a�GB7E�9c�]�K�h��j�iH���>)T�]�q:�n5B,f�(K'��Z�J�9'�赙�!����~�mxV���QK�d���y�x�Sa%����4t4��4[�G�	g��u�ΐ�<�?rd���m�aqw<A�'�����x�]��T���D�սہ��(��I# cg�wr���^���J��VسK���ԝ��y�+M����J۠���� �g��p��Ҩy��\�S>�ī�*:y�g�t?�X)N��8���+�'>_�x'{�g_���ҭ����vb3^���j5CcomO�t�Le�����x��d�a�������}�tS�#BRh��&����<S��݄Ry,����Z&���F
8�琻���G��>S��W��,}7WиWSs��?I���j���2��w����rnKh�3,��\9�צ��Uv��7�x���y�ʂ|v ��m�IY���g}���0�f� r%��Bb^<�K�E�[y�J'K��t��9����~U'#"�>vB�tP,�Q�)6��ߌ�)��3��qL�D �-���x�{��R����Qg{��2�F������=�t1�[)o��ՈPg�Z�����:s/��4A.��N���7�[9_w���-M[��;ZOr��!�Dr�e��u�o�p�>���-��n�m���4����Z��ٛJ���'�1+JH�kh�z�J�G���)f�~��w��&'P�K��Vd�3{�q�u��2��8/���W�I��/[o%]Oa�?Ic-����[Ef6n����%	_��ہ�MA���h�!Vf�݁�/Y��Nռ�Z��8F)"ġ�(���"���ڭ>v��N�?1d�w0���t���Bz�C�m������x����V�$����M{o�=��;d
sJM*��q|����u`f%}�t5��4�����k�xl����f�3_�<�U·���4�����fV�$�C�ʣ"�A�=���$Y	{�d,zs7��)&q̒䔭K.D��C}�G����]F���x�T4��_��u��L�1��0�@$ Oݳ��'��C�H�{���N �'�c�
�˙VC�	n�4�%&B��X�1ucXW�(퓪��M�qZ�����S���N��D��Ӝm@���q�����]{�?O�I��8k���,�'űЮ!%K���S[�cGm�Bl�i��Fؿ�-%6g�ʉ��������=�����!��6x،�{��m}8J��'�Ce��8H ������ҰHOυͰ�rP7�Z�5��$(|�f`ƖYF��]OAa�1���,Y�xc�Q�ê��;u�Ul� �}�H׸�hmO�R�6�i;Bo{QUcחz�^`z�m��tC�+�c\Pʈ���W��1��}t�����.;#:��>�{�l`M�HԠC_��X�En���r�&v��߭֏ܲ��3W��B��B�@7͆y��q96o�+0��q�e��ٙ�`�Q��PК�8Q��_G�����M��~\^:W�Kpe��'�f��1Hf��8Qƿ��
{o��y���uCQ�5�Ȼ�)ȩ�1k�i���ʦ�.�W�oOD[����9�Y�|�Dn���Tk��T�^ZI�>�Z�n��sg�'�)
��?Ҫ�5Wwa5{ޘ�Y�'�4-��� �����w.`+REm�x��h�YsH�����W)�[&��#.\	��5�?�0u�a��;�7�0&Ԥ����jĺ�V+�7>�lM�
[��#l��ʠ�P��b�( g�.��13���Z�R��m��WN�B���\��4�"`��u�=��Đ�N����϶+E�7�i{�����x�|�:�&����H�G�R�U �7[P�j�J����3�1C9`>s�����eo��L���~[�> ުƚ{���8�8�V�L ��3q� 
(��/�9t~��{8j5�I��.����@����j�M�f��f����,S~�R�����컹�� �P�Q�[�t�I��;����i��lʨ��-��S��͂*?�8*U�z�gj���q��o�{*(�hF{A�͠e\�.�<v�ʙ�lKJ�������K�׿�ND��A�zc���#"e��쮌���t֬�S�3�G�] �D2���OY��������EaPz	��U��4��{D����U�82��w~L��P�à��G�0�N젼��r��,���惮r0�!Ak,X��9��6�bv:�����E*6�G���h;����D9���̴�P���-�!��a$�}��`�(w��碡���*�7c,�=�_t��
�� /�h��I~��l(佪�gD䘊��
(�/���	h��~Tǿ��گ�"tk�_9m�� :2�pe_Vgi��P�}�sN��4���i�n0b�_�x���ǜ����5�]���p~���k��1u���s�
r���
�9~̿��u^7��C9�yl6n49S��}����4	�)�Ope2���Q�7�[���=�h��+1[K�žl|�:��a��qbU�qui��m�	93��8xr�Q�7�l���"퍯�YNI�� ��  r�#'/��ݶM���s�Fy~f l���G�����T�(� g�g����k����OB.�}}b��w����<�m�]���Vxk�������楛oZ�����AB����0�X��`���x])0�X��-?�Xy_"@��&z� ���w�'5F��;�uo�7	k.�0�h.��U5�ݢ��_��k�Ě7������i��otYc�/���Q�pכ�ã�`Յ�l�Q��%��q�Bhl�
���ˑT�\&X_�T
�`��ޕ� �p�a	����i��%����_���:�����$�B���^�g�Q�tsW㿅��D�Q��լP�\)�HfX��*	��5�X�4�  `!�!��)�B`_\G(l�] S��5��+	�